// this should be correct
`timescale 1 ns / 1 ns

module testbench();
  logic [13:0] filt_in;
  logic [34:0] filt_out [15:0];
  logic clock, reset, clk_enable;
  logic [13:0] filter_in_data[0:3904];
   
  total_filter filt(.clock(clock), .clk_enable(clk_enable), .reset(reset), .filter_in(filt_in), .filter_out(filt_out));

	always begin
    // clock is correct
		#520;
		clock=~clock;
	end

	initial begin
    clock = 0;
    reset = 1;

    // Input data for filter_in_data_log
    //filter_in_data[0] <= 10'h000;
    //for (int i=1; i<119; i=i+1) filter_in_data[i] <= 10'h200;
    //for (int i=119; i<238; i=i+1) filter_in_data[i] <= 10'h000;
  filter_in_data[   0] <= 14'h1fff;
  filter_in_data[   1] <= 14'h0000;
  filter_in_data[   2] <= 14'h0000;
  filter_in_data[   3] <= 14'h0000;
  filter_in_data[   4] <= 14'h0000;
  filter_in_data[   5] <= 14'h0000;
  filter_in_data[   6] <= 14'h0000;
  filter_in_data[   7] <= 14'h0000;
  filter_in_data[   8] <= 14'h0000;
  filter_in_data[   9] <= 14'h0000;
  filter_in_data[  10] <= 14'h0000;
  filter_in_data[  11] <= 14'h0000;
  filter_in_data[  12] <= 14'h0000;
  filter_in_data[  13] <= 14'h0000;
  filter_in_data[  14] <= 14'h0000;
  filter_in_data[  15] <= 14'h0000;
  filter_in_data[  16] <= 14'h0000;
  filter_in_data[  17] <= 14'h0000;
  filter_in_data[  18] <= 14'h0000;
  filter_in_data[  19] <= 14'h0000;
  filter_in_data[  20] <= 14'h0000;
  filter_in_data[  21] <= 14'h0000;
  filter_in_data[  22] <= 14'h0000;
  filter_in_data[  23] <= 14'h0000;
  filter_in_data[  24] <= 14'h0000;
  filter_in_data[  25] <= 14'h0000;
  filter_in_data[  26] <= 14'h0000;
  filter_in_data[  27] <= 14'h0000;
  filter_in_data[  28] <= 14'h0000;
  filter_in_data[  29] <= 14'h0000;
  filter_in_data[  30] <= 14'h0000;
  filter_in_data[  31] <= 14'h0000;
  filter_in_data[  32] <= 14'h0000;
  filter_in_data[  33] <= 14'h0000;
  filter_in_data[  34] <= 14'h0000;
  filter_in_data[  35] <= 14'h0000;
  filter_in_data[  36] <= 14'h0000;
  filter_in_data[  37] <= 14'h0000;
  filter_in_data[  38] <= 14'h0000;
  filter_in_data[  39] <= 14'h0000;
  filter_in_data[  40] <= 14'h0000;
  filter_in_data[  41] <= 14'h0000;
  filter_in_data[  42] <= 14'h0000;
  filter_in_data[  43] <= 14'h0000;
  filter_in_data[  44] <= 14'h0000;
  filter_in_data[  45] <= 14'h0000;
  filter_in_data[  46] <= 14'h0000;
  filter_in_data[  47] <= 14'h0000;
  filter_in_data[  48] <= 14'h0000;
  filter_in_data[  49] <= 14'h0000;
  filter_in_data[  50] <= 14'h0000;
  filter_in_data[  51] <= 14'h0000;
  filter_in_data[  52] <= 14'h0000;
  filter_in_data[  53] <= 14'h0000;
  filter_in_data[  54] <= 14'h0000;
  filter_in_data[  55] <= 14'h0000;
  filter_in_data[  56] <= 14'h0000;
  filter_in_data[  57] <= 14'h0000;
  filter_in_data[  58] <= 14'h0000;
  filter_in_data[  59] <= 14'h0000;
  filter_in_data[  60] <= 14'h0000;
  filter_in_data[  61] <= 14'h0000;
  filter_in_data[  62] <= 14'h0000;
  filter_in_data[  63] <= 14'h0000;
  filter_in_data[  64] <= 14'h0000;
  filter_in_data[  65] <= 14'h0000;
  filter_in_data[  66] <= 14'h0000;
  filter_in_data[  67] <= 14'h0000;
  filter_in_data[  68] <= 14'h0000;
  filter_in_data[  69] <= 14'h0000;
  filter_in_data[  70] <= 14'h0000;
  filter_in_data[  71] <= 14'h0000;
  filter_in_data[  72] <= 14'h0000;
  filter_in_data[  73] <= 14'h0000;
  filter_in_data[  74] <= 14'h0000;
  filter_in_data[  75] <= 14'h0000;
  filter_in_data[  76] <= 14'h0000;
  filter_in_data[  77] <= 14'h0000;
  filter_in_data[  78] <= 14'h0000;
  filter_in_data[  79] <= 14'h0000;
  filter_in_data[  80] <= 14'h0000;
  filter_in_data[  81] <= 14'h0000;
  filter_in_data[  82] <= 14'h0000;
  filter_in_data[  83] <= 14'h0000;
  filter_in_data[  84] <= 14'h0000;
  filter_in_data[  85] <= 14'h0000;
  filter_in_data[  86] <= 14'h0000;
  filter_in_data[  87] <= 14'h0000;
  filter_in_data[  88] <= 14'h0000;
  filter_in_data[  89] <= 14'h0000;
  filter_in_data[  90] <= 14'h0000;
  filter_in_data[  91] <= 14'h0000;
  filter_in_data[  92] <= 14'h0000;
  filter_in_data[  93] <= 14'h0000;
  filter_in_data[  94] <= 14'h0000;
  filter_in_data[  95] <= 14'h0000;
  filter_in_data[  96] <= 14'h0000;
  filter_in_data[  97] <= 14'h0000;
  filter_in_data[  98] <= 14'h0000;
  filter_in_data[  99] <= 14'h0000;
  filter_in_data[ 100] <= 14'h0000;
  filter_in_data[ 101] <= 14'h0000;
  filter_in_data[ 102] <= 14'h0000;
  filter_in_data[ 103] <= 14'h0000;
  filter_in_data[ 104] <= 14'h0000;
  filter_in_data[ 105] <= 14'h0000;
  filter_in_data[ 106] <= 14'h0000;
  filter_in_data[ 107] <= 14'h0000;
  filter_in_data[ 108] <= 14'h0000;
  filter_in_data[ 109] <= 14'h0000;
  filter_in_data[ 110] <= 14'h0000;
  filter_in_data[ 111] <= 14'h0000;
  filter_in_data[ 112] <= 14'h0000;
  filter_in_data[ 113] <= 14'h0000;
  filter_in_data[ 114] <= 14'h0000;
  filter_in_data[ 115] <= 14'h0000;
  filter_in_data[ 116] <= 14'h0000;
  filter_in_data[ 117] <= 14'h0000;
  filter_in_data[ 118] <= 14'h0000;
  filter_in_data[ 119] <= 14'h0000;
  filter_in_data[ 120] <= 14'h0000;
  filter_in_data[ 121] <= 14'h0000;
  filter_in_data[ 122] <= 14'h0000;
  filter_in_data[ 123] <= 14'h0000;
  filter_in_data[ 124] <= 14'h0000;
  filter_in_data[ 125] <= 14'h0000;
  filter_in_data[ 126] <= 14'h0000;
  filter_in_data[ 127] <= 14'h0000;
  filter_in_data[ 128] <= 14'h0000;
  filter_in_data[ 129] <= 14'h0000;
  filter_in_data[ 130] <= 14'h0000;
  filter_in_data[ 131] <= 14'h0000;
  filter_in_data[ 132] <= 14'h0000;
  filter_in_data[ 133] <= 14'h0000;
  filter_in_data[ 134] <= 14'h0000;
  filter_in_data[ 135] <= 14'h0000;
  filter_in_data[ 136] <= 14'h0000;
  filter_in_data[ 137] <= 14'h0000;
  filter_in_data[ 138] <= 14'h0000;
  filter_in_data[ 139] <= 14'h0000;
  filter_in_data[ 140] <= 14'h0000;
  filter_in_data[ 141] <= 14'h0000;
  filter_in_data[ 142] <= 14'h0000;
  filter_in_data[ 143] <= 14'h0000;
  filter_in_data[ 144] <= 14'h0000;
  filter_in_data[ 145] <= 14'h0000;
  filter_in_data[ 146] <= 14'h0000;
  filter_in_data[ 147] <= 14'h0000;
  filter_in_data[ 148] <= 14'h0000;
  filter_in_data[ 149] <= 14'h0000;
  filter_in_data[ 150] <= 14'h0000;
  filter_in_data[ 151] <= 14'h0000;
  filter_in_data[ 152] <= 14'h0000;
  filter_in_data[ 153] <= 14'h0000;
  filter_in_data[ 154] <= 14'h0000;
  filter_in_data[ 155] <= 14'h0000;
  filter_in_data[ 156] <= 14'h0000;
  filter_in_data[ 157] <= 14'h0000;
  filter_in_data[ 158] <= 14'h0000;
  filter_in_data[ 159] <= 14'h0000;
  filter_in_data[ 160] <= 14'h0000;
  filter_in_data[ 161] <= 14'h0000;
  filter_in_data[ 162] <= 14'h0000;
  filter_in_data[ 163] <= 14'h0000;
  filter_in_data[ 164] <= 14'h0000;
  filter_in_data[ 165] <= 14'h0000;
  filter_in_data[ 166] <= 14'h0000;
  filter_in_data[ 167] <= 14'h0000;
  filter_in_data[ 168] <= 14'h0000;
  filter_in_data[ 169] <= 14'h0000;
  filter_in_data[ 170] <= 14'h0000;
  filter_in_data[ 171] <= 14'h0000;
  filter_in_data[ 172] <= 14'h0000;
  filter_in_data[ 173] <= 14'h0000;
  filter_in_data[ 174] <= 14'h0000;
  filter_in_data[ 175] <= 14'h0000;
  filter_in_data[ 176] <= 14'h0000;
  filter_in_data[ 177] <= 14'h0000;
  filter_in_data[ 178] <= 14'h0000;
  filter_in_data[ 179] <= 14'h0000;
  filter_in_data[ 180] <= 14'h0000;
  filter_in_data[ 181] <= 14'h0000;
  filter_in_data[ 182] <= 14'h0000;
  filter_in_data[ 183] <= 14'h0000;
  filter_in_data[ 184] <= 14'h0000;
  filter_in_data[ 185] <= 14'h0000;
  filter_in_data[ 186] <= 14'h0000;
  filter_in_data[ 187] <= 14'h0000;
  filter_in_data[ 188] <= 14'h0000;
  filter_in_data[ 189] <= 14'h0000;
  filter_in_data[ 190] <= 14'h0000;
  filter_in_data[ 191] <= 14'h0000;
  filter_in_data[ 192] <= 14'h0000;
  filter_in_data[ 193] <= 14'h0000;
  filter_in_data[ 194] <= 14'h0000;
  filter_in_data[ 195] <= 14'h0000;
  filter_in_data[ 196] <= 14'h0000;
  filter_in_data[ 197] <= 14'h0000;
  filter_in_data[ 198] <= 14'h0000;
  filter_in_data[ 199] <= 14'h0000;
  filter_in_data[ 200] <= 14'h0000;
  filter_in_data[ 201] <= 14'h0000;
  filter_in_data[ 202] <= 14'h0000;
  filter_in_data[ 203] <= 14'h0000;
  filter_in_data[ 204] <= 14'h0000;
  filter_in_data[ 205] <= 14'h0000;
  filter_in_data[ 206] <= 14'h0000;
  filter_in_data[ 207] <= 14'h0000;
  filter_in_data[ 208] <= 14'h0000;
  filter_in_data[ 209] <= 14'h0000;
  filter_in_data[ 210] <= 14'h0000;
  filter_in_data[ 211] <= 14'h0000;
  filter_in_data[ 212] <= 14'h0000;
  filter_in_data[ 213] <= 14'h0000;
  filter_in_data[ 214] <= 14'h0000;
  filter_in_data[ 215] <= 14'h0000;
  filter_in_data[ 216] <= 14'h0000;
  filter_in_data[ 217] <= 14'h0000;
  filter_in_data[ 218] <= 14'h0000;
  filter_in_data[ 219] <= 14'h0000;
  filter_in_data[ 220] <= 14'h0000;
  filter_in_data[ 221] <= 14'h0000;
  filter_in_data[ 222] <= 14'h0000;
  filter_in_data[ 223] <= 14'h0000;
  filter_in_data[ 224] <= 14'h0000;
  filter_in_data[ 225] <= 14'h0000;
  filter_in_data[ 226] <= 14'h0000;
  filter_in_data[ 227] <= 14'h0000;
  filter_in_data[ 228] <= 14'h0000;
  filter_in_data[ 229] <= 14'h0000;
  filter_in_data[ 230] <= 14'h0000;
  filter_in_data[ 231] <= 14'h0000;
  filter_in_data[ 232] <= 14'h0000;
  filter_in_data[ 233] <= 14'h0000;
  filter_in_data[ 234] <= 14'h0000;
  filter_in_data[ 235] <= 14'h0000;
  filter_in_data[ 236] <= 14'h0000;
  filter_in_data[ 237] <= 14'h0000;
  filter_in_data[ 238] <= 14'h0000;
  filter_in_data[ 239] <= 14'h1fff;
  filter_in_data[ 240] <= 14'h1fff;
  filter_in_data[ 241] <= 14'h1fff;
  filter_in_data[ 242] <= 14'h1fff;
  filter_in_data[ 243] <= 14'h1fff;
  filter_in_data[ 244] <= 14'h1fff;
  filter_in_data[ 245] <= 14'h1fff;
  filter_in_data[ 246] <= 14'h1fff;
  filter_in_data[ 247] <= 14'h1fff;
  filter_in_data[ 248] <= 14'h1fff;
  filter_in_data[ 249] <= 14'h1fff;
  filter_in_data[ 250] <= 14'h1fff;
  filter_in_data[ 251] <= 14'h1fff;
  filter_in_data[ 252] <= 14'h1fff;
  filter_in_data[ 253] <= 14'h1fff;
  filter_in_data[ 254] <= 14'h1fff;
  filter_in_data[ 255] <= 14'h1fff;
  filter_in_data[ 256] <= 14'h1fff;
  filter_in_data[ 257] <= 14'h1fff;
  filter_in_data[ 258] <= 14'h1fff;
  filter_in_data[ 259] <= 14'h1fff;
  filter_in_data[ 260] <= 14'h1fff;
  filter_in_data[ 261] <= 14'h1fff;
  filter_in_data[ 262] <= 14'h1fff;
  filter_in_data[ 263] <= 14'h1fff;
  filter_in_data[ 264] <= 14'h1fff;
  filter_in_data[ 265] <= 14'h1fff;
  filter_in_data[ 266] <= 14'h1fff;
  filter_in_data[ 267] <= 14'h1fff;
  filter_in_data[ 268] <= 14'h1fff;
  filter_in_data[ 269] <= 14'h1fff;
  filter_in_data[ 270] <= 14'h1fff;
  filter_in_data[ 271] <= 14'h1fff;
  filter_in_data[ 272] <= 14'h1fff;
  filter_in_data[ 273] <= 14'h1fff;
  filter_in_data[ 274] <= 14'h1fff;
  filter_in_data[ 275] <= 14'h1fff;
  filter_in_data[ 276] <= 14'h1fff;
  filter_in_data[ 277] <= 14'h1fff;
  filter_in_data[ 278] <= 14'h1fff;
  filter_in_data[ 279] <= 14'h1fff;
  filter_in_data[ 280] <= 14'h1fff;
  filter_in_data[ 281] <= 14'h1fff;
  filter_in_data[ 282] <= 14'h1fff;
  filter_in_data[ 283] <= 14'h1fff;
  filter_in_data[ 284] <= 14'h1fff;
  filter_in_data[ 285] <= 14'h1fff;
  filter_in_data[ 286] <= 14'h1fff;
  filter_in_data[ 287] <= 14'h1fff;
  filter_in_data[ 288] <= 14'h1fff;
  filter_in_data[ 289] <= 14'h1fff;
  filter_in_data[ 290] <= 14'h1fff;
  filter_in_data[ 291] <= 14'h1fff;
  filter_in_data[ 292] <= 14'h1fff;
  filter_in_data[ 293] <= 14'h1fff;
  filter_in_data[ 294] <= 14'h1fff;
  filter_in_data[ 295] <= 14'h1fff;
  filter_in_data[ 296] <= 14'h1fff;
  filter_in_data[ 297] <= 14'h1fff;
  filter_in_data[ 298] <= 14'h1fff;
  filter_in_data[ 299] <= 14'h1fff;
  filter_in_data[ 300] <= 14'h1fff;
  filter_in_data[ 301] <= 14'h1fff;
  filter_in_data[ 302] <= 14'h1fff;
  filter_in_data[ 303] <= 14'h1fff;
  filter_in_data[ 304] <= 14'h1fff;
  filter_in_data[ 305] <= 14'h1fff;
  filter_in_data[ 306] <= 14'h1fff;
  filter_in_data[ 307] <= 14'h1fff;
  filter_in_data[ 308] <= 14'h1fff;
  filter_in_data[ 309] <= 14'h1fff;
  filter_in_data[ 310] <= 14'h1fff;
  filter_in_data[ 311] <= 14'h1fff;
  filter_in_data[ 312] <= 14'h1fff;
  filter_in_data[ 313] <= 14'h1fff;
  filter_in_data[ 314] <= 14'h1fff;
  filter_in_data[ 315] <= 14'h1fff;
  filter_in_data[ 316] <= 14'h1fff;
  filter_in_data[ 317] <= 14'h1fff;
  filter_in_data[ 318] <= 14'h1fff;
  filter_in_data[ 319] <= 14'h1fff;
  filter_in_data[ 320] <= 14'h1fff;
  filter_in_data[ 321] <= 14'h1fff;
  filter_in_data[ 322] <= 14'h1fff;
  filter_in_data[ 323] <= 14'h1fff;
  filter_in_data[ 324] <= 14'h1fff;
  filter_in_data[ 325] <= 14'h1fff;
  filter_in_data[ 326] <= 14'h1fff;
  filter_in_data[ 327] <= 14'h1fff;
  filter_in_data[ 328] <= 14'h1fff;
  filter_in_data[ 329] <= 14'h1fff;
  filter_in_data[ 330] <= 14'h1fff;
  filter_in_data[ 331] <= 14'h1fff;
  filter_in_data[ 332] <= 14'h1fff;
  filter_in_data[ 333] <= 14'h1fff;
  filter_in_data[ 334] <= 14'h1fff;
  filter_in_data[ 335] <= 14'h1fff;
  filter_in_data[ 336] <= 14'h1fff;
  filter_in_data[ 337] <= 14'h1fff;
  filter_in_data[ 338] <= 14'h1fff;
  filter_in_data[ 339] <= 14'h1fff;
  filter_in_data[ 340] <= 14'h1fff;
  filter_in_data[ 341] <= 14'h1fff;
  filter_in_data[ 342] <= 14'h1fff;
  filter_in_data[ 343] <= 14'h1fff;
  filter_in_data[ 344] <= 14'h1fff;
  filter_in_data[ 345] <= 14'h1fff;
  filter_in_data[ 346] <= 14'h1fff;
  filter_in_data[ 347] <= 14'h1fff;
  filter_in_data[ 348] <= 14'h1fff;
  filter_in_data[ 349] <= 14'h1fff;
  filter_in_data[ 350] <= 14'h1fff;
  filter_in_data[ 351] <= 14'h1fff;
  filter_in_data[ 352] <= 14'h1fff;
  filter_in_data[ 353] <= 14'h1fff;
  filter_in_data[ 354] <= 14'h1fff;
  filter_in_data[ 355] <= 14'h1fff;
  filter_in_data[ 356] <= 14'h1fff;
  filter_in_data[ 357] <= 14'h0000;
  filter_in_data[ 358] <= 14'h0000;
  filter_in_data[ 359] <= 14'h0000;
  filter_in_data[ 360] <= 14'h0000;
  filter_in_data[ 361] <= 14'h0000;
  filter_in_data[ 362] <= 14'h0000;
  filter_in_data[ 363] <= 14'h0000;
  filter_in_data[ 364] <= 14'h0000;
  filter_in_data[ 365] <= 14'h0000;
  filter_in_data[ 366] <= 14'h0000;
  filter_in_data[ 367] <= 14'h0000;
  filter_in_data[ 368] <= 14'h0000;
  filter_in_data[ 369] <= 14'h0000;
  filter_in_data[ 370] <= 14'h0000;
  filter_in_data[ 371] <= 14'h0000;
  filter_in_data[ 372] <= 14'h0000;
  filter_in_data[ 373] <= 14'h0000;
  filter_in_data[ 374] <= 14'h0000;
  filter_in_data[ 375] <= 14'h0000;
  filter_in_data[ 376] <= 14'h0000;
  filter_in_data[ 377] <= 14'h0000;
  filter_in_data[ 378] <= 14'h0000;
  filter_in_data[ 379] <= 14'h0000;
  filter_in_data[ 380] <= 14'h0000;
  filter_in_data[ 381] <= 14'h0000;
  filter_in_data[ 382] <= 14'h0000;
  filter_in_data[ 383] <= 14'h0000;
  filter_in_data[ 384] <= 14'h0000;
  filter_in_data[ 385] <= 14'h0000;
  filter_in_data[ 386] <= 14'h0000;
  filter_in_data[ 387] <= 14'h0000;
  filter_in_data[ 388] <= 14'h0000;
  filter_in_data[ 389] <= 14'h0000;
  filter_in_data[ 390] <= 14'h0000;
  filter_in_data[ 391] <= 14'h0000;
  filter_in_data[ 392] <= 14'h0000;
  filter_in_data[ 393] <= 14'h0000;
  filter_in_data[ 394] <= 14'h0000;
  filter_in_data[ 395] <= 14'h0000;
  filter_in_data[ 396] <= 14'h0000;
  filter_in_data[ 397] <= 14'h0000;
  filter_in_data[ 398] <= 14'h0000;
  filter_in_data[ 399] <= 14'h0000;
  filter_in_data[ 400] <= 14'h0000;
  filter_in_data[ 401] <= 14'h0000;
  filter_in_data[ 402] <= 14'h0000;
  filter_in_data[ 403] <= 14'h0000;
  filter_in_data[ 404] <= 14'h0000;
  filter_in_data[ 405] <= 14'h0000;
  filter_in_data[ 406] <= 14'h0000;
  filter_in_data[ 407] <= 14'h0000;
  filter_in_data[ 408] <= 14'h0000;
  filter_in_data[ 409] <= 14'h0000;
  filter_in_data[ 410] <= 14'h0000;
  filter_in_data[ 411] <= 14'h0000;
  filter_in_data[ 412] <= 14'h0000;
  filter_in_data[ 413] <= 14'h0000;
  filter_in_data[ 414] <= 14'h0000;
  filter_in_data[ 415] <= 14'h0000;
  filter_in_data[ 416] <= 14'h0000;
  filter_in_data[ 417] <= 14'h0000;
  filter_in_data[ 418] <= 14'h0000;
  filter_in_data[ 419] <= 14'h0000;
  filter_in_data[ 420] <= 14'h0000;
  filter_in_data[ 421] <= 14'h0000;
  filter_in_data[ 422] <= 14'h0000;
  filter_in_data[ 423] <= 14'h0000;
  filter_in_data[ 424] <= 14'h0000;
  filter_in_data[ 425] <= 14'h0000;
  filter_in_data[ 426] <= 14'h0000;
  filter_in_data[ 427] <= 14'h0000;
  filter_in_data[ 428] <= 14'h0000;
  filter_in_data[ 429] <= 14'h0000;
  filter_in_data[ 430] <= 14'h0000;
  filter_in_data[ 431] <= 14'h0000;
  filter_in_data[ 432] <= 14'h0000;
  filter_in_data[ 433] <= 14'h0000;
  filter_in_data[ 434] <= 14'h0000;
  filter_in_data[ 435] <= 14'h0000;
  filter_in_data[ 436] <= 14'h0000;
  filter_in_data[ 437] <= 14'h0000;
  filter_in_data[ 438] <= 14'h0000;
  filter_in_data[ 439] <= 14'h0000;
  filter_in_data[ 440] <= 14'h0000;
  filter_in_data[ 441] <= 14'h0000;
  filter_in_data[ 442] <= 14'h0000;
  filter_in_data[ 443] <= 14'h0000;
  filter_in_data[ 444] <= 14'h0000;
  filter_in_data[ 445] <= 14'h0000;
  filter_in_data[ 446] <= 14'h0000;
  filter_in_data[ 447] <= 14'h0000;
  filter_in_data[ 448] <= 14'h0000;
  filter_in_data[ 449] <= 14'h0000;
  filter_in_data[ 450] <= 14'h0000;
  filter_in_data[ 451] <= 14'h0000;
  filter_in_data[ 452] <= 14'h0000;
  filter_in_data[ 453] <= 14'h0000;
  filter_in_data[ 454] <= 14'h0000;
  filter_in_data[ 455] <= 14'h0000;
  filter_in_data[ 456] <= 14'h0000;
  filter_in_data[ 457] <= 14'h0000;
  filter_in_data[ 458] <= 14'h0000;
  filter_in_data[ 459] <= 14'h0000;
  filter_in_data[ 460] <= 14'h0000;
  filter_in_data[ 461] <= 14'h0000;
  filter_in_data[ 462] <= 14'h0000;
  filter_in_data[ 463] <= 14'h0000;
  filter_in_data[ 464] <= 14'h0000;
  filter_in_data[ 465] <= 14'h0000;
  filter_in_data[ 466] <= 14'h0000;
  filter_in_data[ 467] <= 14'h0000;
  filter_in_data[ 468] <= 14'h0000;
  filter_in_data[ 469] <= 14'h0000;
  filter_in_data[ 470] <= 14'h0000;
  filter_in_data[ 471] <= 14'h0000;
  filter_in_data[ 472] <= 14'h0000;
  filter_in_data[ 473] <= 14'h0000;
  filter_in_data[ 474] <= 14'h0000;
  filter_in_data[ 475] <= 14'h0000;
  filter_in_data[ 476] <= 14'h2000;
  filter_in_data[ 477] <= 14'h2010;
  filter_in_data[ 478] <= 14'h2020;
  filter_in_data[ 479] <= 14'h2030;
  filter_in_data[ 480] <= 14'h2040;
  filter_in_data[ 481] <= 14'h2050;
  filter_in_data[ 482] <= 14'h2060;
  filter_in_data[ 483] <= 14'h2070;
  filter_in_data[ 484] <= 14'h2080;
  filter_in_data[ 485] <= 14'h2090;
  filter_in_data[ 486] <= 14'h20a0;
  filter_in_data[ 487] <= 14'h20b0;
  filter_in_data[ 488] <= 14'h20c0;
  filter_in_data[ 489] <= 14'h20d0;
  filter_in_data[ 490] <= 14'h20e0;
  filter_in_data[ 491] <= 14'h20f0;
  filter_in_data[ 492] <= 14'h2100;
  filter_in_data[ 493] <= 14'h2110;
  filter_in_data[ 494] <= 14'h2120;
  filter_in_data[ 495] <= 14'h2130;
  filter_in_data[ 496] <= 14'h2140;
  filter_in_data[ 497] <= 14'h2150;
  filter_in_data[ 498] <= 14'h2160;
  filter_in_data[ 499] <= 14'h2170;
  filter_in_data[ 500] <= 14'h2180;
  filter_in_data[ 501] <= 14'h2190;
  filter_in_data[ 502] <= 14'h21a0;
  filter_in_data[ 503] <= 14'h21b0;
  filter_in_data[ 504] <= 14'h21c0;
  filter_in_data[ 505] <= 14'h21d0;
  filter_in_data[ 506] <= 14'h21e0;
  filter_in_data[ 507] <= 14'h21f0;
  filter_in_data[ 508] <= 14'h2201;
  filter_in_data[ 509] <= 14'h2211;
  filter_in_data[ 510] <= 14'h2221;
  filter_in_data[ 511] <= 14'h2231;
  filter_in_data[ 512] <= 14'h2241;
  filter_in_data[ 513] <= 14'h2251;
  filter_in_data[ 514] <= 14'h2261;
  filter_in_data[ 515] <= 14'h2271;
  filter_in_data[ 516] <= 14'h2281;
  filter_in_data[ 517] <= 14'h2291;
  filter_in_data[ 518] <= 14'h22a1;
  filter_in_data[ 519] <= 14'h22b1;
  filter_in_data[ 520] <= 14'h22c1;
  filter_in_data[ 521] <= 14'h22d1;
  filter_in_data[ 522] <= 14'h22e1;
  filter_in_data[ 523] <= 14'h22f1;
  filter_in_data[ 524] <= 14'h2301;
  filter_in_data[ 525] <= 14'h2311;
  filter_in_data[ 526] <= 14'h2321;
  filter_in_data[ 527] <= 14'h2331;
  filter_in_data[ 528] <= 14'h2341;
  filter_in_data[ 529] <= 14'h2351;
  filter_in_data[ 530] <= 14'h2361;
  filter_in_data[ 531] <= 14'h2371;
  filter_in_data[ 532] <= 14'h2381;
  filter_in_data[ 533] <= 14'h2391;
  filter_in_data[ 534] <= 14'h23a1;
  filter_in_data[ 535] <= 14'h23b1;
  filter_in_data[ 536] <= 14'h23c1;
  filter_in_data[ 537] <= 14'h23d1;
  filter_in_data[ 538] <= 14'h23e1;
  filter_in_data[ 539] <= 14'h23f1;
  filter_in_data[ 540] <= 14'h2401;
  filter_in_data[ 541] <= 14'h2411;
  filter_in_data[ 542] <= 14'h2421;
  filter_in_data[ 543] <= 14'h2431;
  filter_in_data[ 544] <= 14'h2441;
  filter_in_data[ 545] <= 14'h2451;
  filter_in_data[ 546] <= 14'h2461;
  filter_in_data[ 547] <= 14'h2471;
  filter_in_data[ 548] <= 14'h2481;
  filter_in_data[ 549] <= 14'h2491;
  filter_in_data[ 550] <= 14'h24a1;
  filter_in_data[ 551] <= 14'h24b1;
  filter_in_data[ 552] <= 14'h24c1;
  filter_in_data[ 553] <= 14'h24d1;
  filter_in_data[ 554] <= 14'h24e1;
  filter_in_data[ 555] <= 14'h24f1;
  filter_in_data[ 556] <= 14'h2501;
  filter_in_data[ 557] <= 14'h2511;
  filter_in_data[ 558] <= 14'h2521;
  filter_in_data[ 559] <= 14'h2531;
  filter_in_data[ 560] <= 14'h2541;
  filter_in_data[ 561] <= 14'h2551;
  filter_in_data[ 562] <= 14'h2561;
  filter_in_data[ 563] <= 14'h2571;
  filter_in_data[ 564] <= 14'h2581;
  filter_in_data[ 565] <= 14'h2591;
  filter_in_data[ 566] <= 14'h25a1;
  filter_in_data[ 567] <= 14'h25b1;
  filter_in_data[ 568] <= 14'h25c1;
  filter_in_data[ 569] <= 14'h25d1;
  filter_in_data[ 570] <= 14'h25e1;
  filter_in_data[ 571] <= 14'h25f1;
  filter_in_data[ 572] <= 14'h2602;
  filter_in_data[ 573] <= 14'h2612;
  filter_in_data[ 574] <= 14'h2622;
  filter_in_data[ 575] <= 14'h2632;
  filter_in_data[ 576] <= 14'h2642;
  filter_in_data[ 577] <= 14'h2652;
  filter_in_data[ 578] <= 14'h2662;
  filter_in_data[ 579] <= 14'h2672;
  filter_in_data[ 580] <= 14'h2682;
  filter_in_data[ 581] <= 14'h2692;
  filter_in_data[ 582] <= 14'h26a2;
  filter_in_data[ 583] <= 14'h26b2;
  filter_in_data[ 584] <= 14'h26c2;
  filter_in_data[ 585] <= 14'h26d2;
  filter_in_data[ 586] <= 14'h26e2;
  filter_in_data[ 587] <= 14'h26f2;
  filter_in_data[ 588] <= 14'h2702;
  filter_in_data[ 589] <= 14'h2712;
  filter_in_data[ 590] <= 14'h2722;
  filter_in_data[ 591] <= 14'h2732;
  filter_in_data[ 592] <= 14'h2742;
  filter_in_data[ 593] <= 14'h2752;
  filter_in_data[ 594] <= 14'h2762;
  filter_in_data[ 595] <= 14'h2772;
  filter_in_data[ 596] <= 14'h2782;
  filter_in_data[ 597] <= 14'h2792;
  filter_in_data[ 598] <= 14'h27a2;
  filter_in_data[ 599] <= 14'h27b2;
  filter_in_data[ 600] <= 14'h27c2;
  filter_in_data[ 601] <= 14'h27d2;
  filter_in_data[ 602] <= 14'h27e2;
  filter_in_data[ 603] <= 14'h27f2;
  filter_in_data[ 604] <= 14'h2802;
  filter_in_data[ 605] <= 14'h2812;
  filter_in_data[ 606] <= 14'h2822;
  filter_in_data[ 607] <= 14'h2832;
  filter_in_data[ 608] <= 14'h2842;
  filter_in_data[ 609] <= 14'h2852;
  filter_in_data[ 610] <= 14'h2862;
  filter_in_data[ 611] <= 14'h2872;
  filter_in_data[ 612] <= 14'h2882;
  filter_in_data[ 613] <= 14'h2892;
  filter_in_data[ 614] <= 14'h28a2;
  filter_in_data[ 615] <= 14'h28b2;
  filter_in_data[ 616] <= 14'h28c2;
  filter_in_data[ 617] <= 14'h28d2;
  filter_in_data[ 618] <= 14'h28e2;
  filter_in_data[ 619] <= 14'h28f2;
  filter_in_data[ 620] <= 14'h2902;
  filter_in_data[ 621] <= 14'h2912;
  filter_in_data[ 622] <= 14'h2922;
  filter_in_data[ 623] <= 14'h2932;
  filter_in_data[ 624] <= 14'h2942;
  filter_in_data[ 625] <= 14'h2952;
  filter_in_data[ 626] <= 14'h2962;
  filter_in_data[ 627] <= 14'h2972;
  filter_in_data[ 628] <= 14'h2982;
  filter_in_data[ 629] <= 14'h2992;
  filter_in_data[ 630] <= 14'h29a2;
  filter_in_data[ 631] <= 14'h29b2;
  filter_in_data[ 632] <= 14'h29c2;
  filter_in_data[ 633] <= 14'h29d2;
  filter_in_data[ 634] <= 14'h29e2;
  filter_in_data[ 635] <= 14'h29f2;
  filter_in_data[ 636] <= 14'h2a03;
  filter_in_data[ 637] <= 14'h2a13;
  filter_in_data[ 638] <= 14'h2a23;
  filter_in_data[ 639] <= 14'h2a33;
  filter_in_data[ 640] <= 14'h2a43;
  filter_in_data[ 641] <= 14'h2a53;
  filter_in_data[ 642] <= 14'h2a63;
  filter_in_data[ 643] <= 14'h2a73;
  filter_in_data[ 644] <= 14'h2a83;
  filter_in_data[ 645] <= 14'h2a93;
  filter_in_data[ 646] <= 14'h2aa3;
  filter_in_data[ 647] <= 14'h2ab3;
  filter_in_data[ 648] <= 14'h2ac3;
  filter_in_data[ 649] <= 14'h2ad3;
  filter_in_data[ 650] <= 14'h2ae3;
  filter_in_data[ 651] <= 14'h2af3;
  filter_in_data[ 652] <= 14'h2b03;
  filter_in_data[ 653] <= 14'h2b13;
  filter_in_data[ 654] <= 14'h2b23;
  filter_in_data[ 655] <= 14'h2b33;
  filter_in_data[ 656] <= 14'h2b43;
  filter_in_data[ 657] <= 14'h2b53;
  filter_in_data[ 658] <= 14'h2b63;
  filter_in_data[ 659] <= 14'h2b73;
  filter_in_data[ 660] <= 14'h2b83;
  filter_in_data[ 661] <= 14'h2b93;
  filter_in_data[ 662] <= 14'h2ba3;
  filter_in_data[ 663] <= 14'h2bb3;
  filter_in_data[ 664] <= 14'h2bc3;
  filter_in_data[ 665] <= 14'h2bd3;
  filter_in_data[ 666] <= 14'h2be3;
  filter_in_data[ 667] <= 14'h2bf3;
  filter_in_data[ 668] <= 14'h2c03;
  filter_in_data[ 669] <= 14'h2c13;
  filter_in_data[ 670] <= 14'h2c23;
  filter_in_data[ 671] <= 14'h2c33;
  filter_in_data[ 672] <= 14'h2c43;
  filter_in_data[ 673] <= 14'h2c53;
  filter_in_data[ 674] <= 14'h2c63;
  filter_in_data[ 675] <= 14'h2c73;
  filter_in_data[ 676] <= 14'h2c83;
  filter_in_data[ 677] <= 14'h2c93;
  filter_in_data[ 678] <= 14'h2ca3;
  filter_in_data[ 679] <= 14'h2cb3;
  filter_in_data[ 680] <= 14'h2cc3;
  filter_in_data[ 681] <= 14'h2cd3;
  filter_in_data[ 682] <= 14'h2ce3;
  filter_in_data[ 683] <= 14'h2cf3;
  filter_in_data[ 684] <= 14'h2d03;
  filter_in_data[ 685] <= 14'h2d13;
  filter_in_data[ 686] <= 14'h2d23;
  filter_in_data[ 687] <= 14'h2d33;
  filter_in_data[ 688] <= 14'h2d43;
  filter_in_data[ 689] <= 14'h2d53;
  filter_in_data[ 690] <= 14'h2d63;
  filter_in_data[ 691] <= 14'h2d73;
  filter_in_data[ 692] <= 14'h2d83;
  filter_in_data[ 693] <= 14'h2d93;
  filter_in_data[ 694] <= 14'h2da3;
  filter_in_data[ 695] <= 14'h2db3;
  filter_in_data[ 696] <= 14'h2dc3;
  filter_in_data[ 697] <= 14'h2dd3;
  filter_in_data[ 698] <= 14'h2de3;
  filter_in_data[ 699] <= 14'h2df3;
  filter_in_data[ 700] <= 14'h2e04;
  filter_in_data[ 701] <= 14'h2e14;
  filter_in_data[ 702] <= 14'h2e24;
  filter_in_data[ 703] <= 14'h2e34;
  filter_in_data[ 704] <= 14'h2e44;
  filter_in_data[ 705] <= 14'h2e54;
  filter_in_data[ 706] <= 14'h2e64;
  filter_in_data[ 707] <= 14'h2e74;
  filter_in_data[ 708] <= 14'h2e84;
  filter_in_data[ 709] <= 14'h2e94;
  filter_in_data[ 710] <= 14'h2ea4;
  filter_in_data[ 711] <= 14'h2eb4;
  filter_in_data[ 712] <= 14'h2ec4;
  filter_in_data[ 713] <= 14'h2ed4;
  filter_in_data[ 714] <= 14'h2ee4;
  filter_in_data[ 715] <= 14'h2ef4;
  filter_in_data[ 716] <= 14'h2f04;
  filter_in_data[ 717] <= 14'h2f14;
  filter_in_data[ 718] <= 14'h2f24;
  filter_in_data[ 719] <= 14'h2f34;
  filter_in_data[ 720] <= 14'h2f44;
  filter_in_data[ 721] <= 14'h2f54;
  filter_in_data[ 722] <= 14'h2f64;
  filter_in_data[ 723] <= 14'h2f74;
  filter_in_data[ 724] <= 14'h2f84;
  filter_in_data[ 725] <= 14'h2f94;
  filter_in_data[ 726] <= 14'h2fa4;
  filter_in_data[ 727] <= 14'h2fb4;
  filter_in_data[ 728] <= 14'h2fc4;
  filter_in_data[ 729] <= 14'h2fd4;
  filter_in_data[ 730] <= 14'h2fe4;
  filter_in_data[ 731] <= 14'h2ff4;
  filter_in_data[ 732] <= 14'h3004;
  filter_in_data[ 733] <= 14'h3014;
  filter_in_data[ 734] <= 14'h3024;
  filter_in_data[ 735] <= 14'h3034;
  filter_in_data[ 736] <= 14'h3044;
  filter_in_data[ 737] <= 14'h3054;
  filter_in_data[ 738] <= 14'h3064;
  filter_in_data[ 739] <= 14'h3074;
  filter_in_data[ 740] <= 14'h3084;
  filter_in_data[ 741] <= 14'h3094;
  filter_in_data[ 742] <= 14'h30a4;
  filter_in_data[ 743] <= 14'h30b4;
  filter_in_data[ 744] <= 14'h30c4;
  filter_in_data[ 745] <= 14'h30d4;
  filter_in_data[ 746] <= 14'h30e4;
  filter_in_data[ 747] <= 14'h30f4;
  filter_in_data[ 748] <= 14'h3104;
  filter_in_data[ 749] <= 14'h3114;
  filter_in_data[ 750] <= 14'h3124;
  filter_in_data[ 751] <= 14'h3134;
  filter_in_data[ 752] <= 14'h3144;
  filter_in_data[ 753] <= 14'h3154;
  filter_in_data[ 754] <= 14'h3164;
  filter_in_data[ 755] <= 14'h3174;
  filter_in_data[ 756] <= 14'h3184;
  filter_in_data[ 757] <= 14'h3194;
  filter_in_data[ 758] <= 14'h31a4;
  filter_in_data[ 759] <= 14'h31b4;
  filter_in_data[ 760] <= 14'h31c4;
  filter_in_data[ 761] <= 14'h31d4;
  filter_in_data[ 762] <= 14'h31e4;
  filter_in_data[ 763] <= 14'h31f4;
  filter_in_data[ 764] <= 14'h3205;
  filter_in_data[ 765] <= 14'h3215;
  filter_in_data[ 766] <= 14'h3225;
  filter_in_data[ 767] <= 14'h3235;
  filter_in_data[ 768] <= 14'h3245;
  filter_in_data[ 769] <= 14'h3255;
  filter_in_data[ 770] <= 14'h3265;
  filter_in_data[ 771] <= 14'h3275;
  filter_in_data[ 772] <= 14'h3285;
  filter_in_data[ 773] <= 14'h3295;
  filter_in_data[ 774] <= 14'h32a5;
  filter_in_data[ 775] <= 14'h32b5;
  filter_in_data[ 776] <= 14'h32c5;
  filter_in_data[ 777] <= 14'h32d5;
  filter_in_data[ 778] <= 14'h32e5;
  filter_in_data[ 779] <= 14'h32f5;
  filter_in_data[ 780] <= 14'h3305;
  filter_in_data[ 781] <= 14'h3315;
  filter_in_data[ 782] <= 14'h3325;
  filter_in_data[ 783] <= 14'h3335;
  filter_in_data[ 784] <= 14'h3345;
  filter_in_data[ 785] <= 14'h3355;
  filter_in_data[ 786] <= 14'h3365;
  filter_in_data[ 787] <= 14'h3375;
  filter_in_data[ 788] <= 14'h3385;
  filter_in_data[ 789] <= 14'h3395;
  filter_in_data[ 790] <= 14'h33a5;
  filter_in_data[ 791] <= 14'h33b5;
  filter_in_data[ 792] <= 14'h33c5;
  filter_in_data[ 793] <= 14'h33d5;
  filter_in_data[ 794] <= 14'h33e5;
  filter_in_data[ 795] <= 14'h33f5;
  filter_in_data[ 796] <= 14'h3405;
  filter_in_data[ 797] <= 14'h3415;
  filter_in_data[ 798] <= 14'h3425;
  filter_in_data[ 799] <= 14'h3435;
  filter_in_data[ 800] <= 14'h3445;
  filter_in_data[ 801] <= 14'h3455;
  filter_in_data[ 802] <= 14'h3465;
  filter_in_data[ 803] <= 14'h3475;
  filter_in_data[ 804] <= 14'h3485;
  filter_in_data[ 805] <= 14'h3495;
  filter_in_data[ 806] <= 14'h34a5;
  filter_in_data[ 807] <= 14'h34b5;
  filter_in_data[ 808] <= 14'h34c5;
  filter_in_data[ 809] <= 14'h34d5;
  filter_in_data[ 810] <= 14'h34e5;
  filter_in_data[ 811] <= 14'h34f5;
  filter_in_data[ 812] <= 14'h3505;
  filter_in_data[ 813] <= 14'h3515;
  filter_in_data[ 814] <= 14'h3525;
  filter_in_data[ 815] <= 14'h3535;
  filter_in_data[ 816] <= 14'h3545;
  filter_in_data[ 817] <= 14'h3555;
  filter_in_data[ 818] <= 14'h3565;
  filter_in_data[ 819] <= 14'h3575;
  filter_in_data[ 820] <= 14'h3585;
  filter_in_data[ 821] <= 14'h3595;
  filter_in_data[ 822] <= 14'h35a5;
  filter_in_data[ 823] <= 14'h35b5;
  filter_in_data[ 824] <= 14'h35c5;
  filter_in_data[ 825] <= 14'h35d5;
  filter_in_data[ 826] <= 14'h35e5;
  filter_in_data[ 827] <= 14'h35f5;
  filter_in_data[ 828] <= 14'h3606;
  filter_in_data[ 829] <= 14'h3616;
  filter_in_data[ 830] <= 14'h3626;
  filter_in_data[ 831] <= 14'h3636;
  filter_in_data[ 832] <= 14'h3646;
  filter_in_data[ 833] <= 14'h3656;
  filter_in_data[ 834] <= 14'h3666;
  filter_in_data[ 835] <= 14'h3676;
  filter_in_data[ 836] <= 14'h3686;
  filter_in_data[ 837] <= 14'h3696;
  filter_in_data[ 838] <= 14'h36a6;
  filter_in_data[ 839] <= 14'h36b6;
  filter_in_data[ 840] <= 14'h36c6;
  filter_in_data[ 841] <= 14'h36d6;
  filter_in_data[ 842] <= 14'h36e6;
  filter_in_data[ 843] <= 14'h36f6;
  filter_in_data[ 844] <= 14'h3706;
  filter_in_data[ 845] <= 14'h3716;
  filter_in_data[ 846] <= 14'h3726;
  filter_in_data[ 847] <= 14'h3736;
  filter_in_data[ 848] <= 14'h3746;
  filter_in_data[ 849] <= 14'h3756;
  filter_in_data[ 850] <= 14'h3766;
  filter_in_data[ 851] <= 14'h3776;
  filter_in_data[ 852] <= 14'h3786;
  filter_in_data[ 853] <= 14'h3796;
  filter_in_data[ 854] <= 14'h37a6;
  filter_in_data[ 855] <= 14'h37b6;
  filter_in_data[ 856] <= 14'h37c6;
  filter_in_data[ 857] <= 14'h37d6;
  filter_in_data[ 858] <= 14'h37e6;
  filter_in_data[ 859] <= 14'h37f6;
  filter_in_data[ 860] <= 14'h3806;
  filter_in_data[ 861] <= 14'h3816;
  filter_in_data[ 862] <= 14'h3826;
  filter_in_data[ 863] <= 14'h3836;
  filter_in_data[ 864] <= 14'h3846;
  filter_in_data[ 865] <= 14'h3856;
  filter_in_data[ 866] <= 14'h3866;
  filter_in_data[ 867] <= 14'h3876;
  filter_in_data[ 868] <= 14'h3886;
  filter_in_data[ 869] <= 14'h3896;
  filter_in_data[ 870] <= 14'h38a6;
  filter_in_data[ 871] <= 14'h38b6;
  filter_in_data[ 872] <= 14'h38c6;
  filter_in_data[ 873] <= 14'h38d6;
  filter_in_data[ 874] <= 14'h38e6;
  filter_in_data[ 875] <= 14'h38f6;
  filter_in_data[ 876] <= 14'h3906;
  filter_in_data[ 877] <= 14'h3916;
  filter_in_data[ 878] <= 14'h3926;
  filter_in_data[ 879] <= 14'h3936;
  filter_in_data[ 880] <= 14'h3946;
  filter_in_data[ 881] <= 14'h3956;
  filter_in_data[ 882] <= 14'h3966;
  filter_in_data[ 883] <= 14'h3976;
  filter_in_data[ 884] <= 14'h3986;
  filter_in_data[ 885] <= 14'h3996;
  filter_in_data[ 886] <= 14'h39a6;
  filter_in_data[ 887] <= 14'h39b6;
  filter_in_data[ 888] <= 14'h39c6;
  filter_in_data[ 889] <= 14'h39d6;
  filter_in_data[ 890] <= 14'h39e6;
  filter_in_data[ 891] <= 14'h39f6;
  filter_in_data[ 892] <= 14'h3a07;
  filter_in_data[ 893] <= 14'h3a17;
  filter_in_data[ 894] <= 14'h3a27;
  filter_in_data[ 895] <= 14'h3a37;
  filter_in_data[ 896] <= 14'h3a47;
  filter_in_data[ 897] <= 14'h3a57;
  filter_in_data[ 898] <= 14'h3a67;
  filter_in_data[ 899] <= 14'h3a77;
  filter_in_data[ 900] <= 14'h3a87;
  filter_in_data[ 901] <= 14'h3a97;
  filter_in_data[ 902] <= 14'h3aa7;
  filter_in_data[ 903] <= 14'h3ab7;
  filter_in_data[ 904] <= 14'h3ac7;
  filter_in_data[ 905] <= 14'h3ad7;
  filter_in_data[ 906] <= 14'h3ae7;
  filter_in_data[ 907] <= 14'h3af7;
  filter_in_data[ 908] <= 14'h3b07;
  filter_in_data[ 909] <= 14'h3b17;
  filter_in_data[ 910] <= 14'h3b27;
  filter_in_data[ 911] <= 14'h3b37;
  filter_in_data[ 912] <= 14'h3b47;
  filter_in_data[ 913] <= 14'h3b57;
  filter_in_data[ 914] <= 14'h3b67;
  filter_in_data[ 915] <= 14'h3b77;
  filter_in_data[ 916] <= 14'h3b87;
  filter_in_data[ 917] <= 14'h3b97;
  filter_in_data[ 918] <= 14'h3ba7;
  filter_in_data[ 919] <= 14'h3bb7;
  filter_in_data[ 920] <= 14'h3bc7;
  filter_in_data[ 921] <= 14'h3bd7;
  filter_in_data[ 922] <= 14'h3be7;
  filter_in_data[ 923] <= 14'h3bf7;
  filter_in_data[ 924] <= 14'h3c07;
  filter_in_data[ 925] <= 14'h3c17;
  filter_in_data[ 926] <= 14'h3c27;
  filter_in_data[ 927] <= 14'h3c37;
  filter_in_data[ 928] <= 14'h3c47;
  filter_in_data[ 929] <= 14'h3c57;
  filter_in_data[ 930] <= 14'h3c67;
  filter_in_data[ 931] <= 14'h3c77;
  filter_in_data[ 932] <= 14'h3c87;
  filter_in_data[ 933] <= 14'h3c97;
  filter_in_data[ 934] <= 14'h3ca7;
  filter_in_data[ 935] <= 14'h3cb7;
  filter_in_data[ 936] <= 14'h3cc7;
  filter_in_data[ 937] <= 14'h3cd7;
  filter_in_data[ 938] <= 14'h3ce7;
  filter_in_data[ 939] <= 14'h3cf7;
  filter_in_data[ 940] <= 14'h3d07;
  filter_in_data[ 941] <= 14'h3d17;
  filter_in_data[ 942] <= 14'h3d27;
  filter_in_data[ 943] <= 14'h3d37;
  filter_in_data[ 944] <= 14'h3d47;
  filter_in_data[ 945] <= 14'h3d57;
  filter_in_data[ 946] <= 14'h3d67;
  filter_in_data[ 947] <= 14'h3d77;
  filter_in_data[ 948] <= 14'h3d87;
  filter_in_data[ 949] <= 14'h3d97;
  filter_in_data[ 950] <= 14'h3da7;
  filter_in_data[ 951] <= 14'h3db7;
  filter_in_data[ 952] <= 14'h3dc7;
  filter_in_data[ 953] <= 14'h3dd7;
  filter_in_data[ 954] <= 14'h3de7;
  filter_in_data[ 955] <= 14'h3df7;
  filter_in_data[ 956] <= 14'h3e08;
  filter_in_data[ 957] <= 14'h3e18;
  filter_in_data[ 958] <= 14'h3e28;
  filter_in_data[ 959] <= 14'h3e38;
  filter_in_data[ 960] <= 14'h3e48;
  filter_in_data[ 961] <= 14'h3e58;
  filter_in_data[ 962] <= 14'h3e68;
  filter_in_data[ 963] <= 14'h3e78;
  filter_in_data[ 964] <= 14'h3e88;
  filter_in_data[ 965] <= 14'h3e98;
  filter_in_data[ 966] <= 14'h3ea8;
  filter_in_data[ 967] <= 14'h3eb8;
  filter_in_data[ 968] <= 14'h3ec8;
  filter_in_data[ 969] <= 14'h3ed8;
  filter_in_data[ 970] <= 14'h3ee8;
  filter_in_data[ 971] <= 14'h3ef8;
  filter_in_data[ 972] <= 14'h3f08;
  filter_in_data[ 973] <= 14'h3f18;
  filter_in_data[ 974] <= 14'h3f28;
  filter_in_data[ 975] <= 14'h3f38;
  filter_in_data[ 976] <= 14'h3f48;
  filter_in_data[ 977] <= 14'h3f58;
  filter_in_data[ 978] <= 14'h3f68;
  filter_in_data[ 979] <= 14'h3f78;
  filter_in_data[ 980] <= 14'h3f88;
  filter_in_data[ 981] <= 14'h3f98;
  filter_in_data[ 982] <= 14'h3fa8;
  filter_in_data[ 983] <= 14'h3fb8;
  filter_in_data[ 984] <= 14'h3fc8;
  filter_in_data[ 985] <= 14'h3fd8;
  filter_in_data[ 986] <= 14'h3fe8;
  filter_in_data[ 987] <= 14'h3ff8;
  filter_in_data[ 988] <= 14'h0008;
  filter_in_data[ 989] <= 14'h0018;
  filter_in_data[ 990] <= 14'h0028;
  filter_in_data[ 991] <= 14'h0038;
  filter_in_data[ 992] <= 14'h0048;
  filter_in_data[ 993] <= 14'h0058;
  filter_in_data[ 994] <= 14'h0068;
  filter_in_data[ 995] <= 14'h0078;
  filter_in_data[ 996] <= 14'h0088;
  filter_in_data[ 997] <= 14'h0098;
  filter_in_data[ 998] <= 14'h00a8;
  filter_in_data[ 999] <= 14'h00b8;
  filter_in_data[1000] <= 14'h00c8;
  filter_in_data[1001] <= 14'h00d8;
  filter_in_data[1002] <= 14'h00e8;
  filter_in_data[1003] <= 14'h00f8;
  filter_in_data[1004] <= 14'h0108;
  filter_in_data[1005] <= 14'h0118;
  filter_in_data[1006] <= 14'h0128;
  filter_in_data[1007] <= 14'h0138;
  filter_in_data[1008] <= 14'h0148;
  filter_in_data[1009] <= 14'h0158;
  filter_in_data[1010] <= 14'h0168;
  filter_in_data[1011] <= 14'h0178;
  filter_in_data[1012] <= 14'h0188;
  filter_in_data[1013] <= 14'h0198;
  filter_in_data[1014] <= 14'h01a8;
  filter_in_data[1015] <= 14'h01b8;
  filter_in_data[1016] <= 14'h01c8;
  filter_in_data[1017] <= 14'h01d8;
  filter_in_data[1018] <= 14'h01e8;
  filter_in_data[1019] <= 14'h01f8;
  filter_in_data[1020] <= 14'h0209;
  filter_in_data[1021] <= 14'h0219;
  filter_in_data[1022] <= 14'h0229;
  filter_in_data[1023] <= 14'h0239;
  filter_in_data[1024] <= 14'h0249;
  filter_in_data[1025] <= 14'h0259;
  filter_in_data[1026] <= 14'h0269;
  filter_in_data[1027] <= 14'h0279;
  filter_in_data[1028] <= 14'h0289;
  filter_in_data[1029] <= 14'h0299;
  filter_in_data[1030] <= 14'h02a9;
  filter_in_data[1031] <= 14'h02b9;
  filter_in_data[1032] <= 14'h02c9;
  filter_in_data[1033] <= 14'h02d9;
  filter_in_data[1034] <= 14'h02e9;
  filter_in_data[1035] <= 14'h02f9;
  filter_in_data[1036] <= 14'h0309;
  filter_in_data[1037] <= 14'h0319;
  filter_in_data[1038] <= 14'h0329;
  filter_in_data[1039] <= 14'h0339;
  filter_in_data[1040] <= 14'h0349;
  filter_in_data[1041] <= 14'h0359;
  filter_in_data[1042] <= 14'h0369;
  filter_in_data[1043] <= 14'h0379;
  filter_in_data[1044] <= 14'h0389;
  filter_in_data[1045] <= 14'h0399;
  filter_in_data[1046] <= 14'h03a9;
  filter_in_data[1047] <= 14'h03b9;
  filter_in_data[1048] <= 14'h03c9;
  filter_in_data[1049] <= 14'h03d9;
  filter_in_data[1050] <= 14'h03e9;
  filter_in_data[1051] <= 14'h03f9;
  filter_in_data[1052] <= 14'h0409;
  filter_in_data[1053] <= 14'h0419;
  filter_in_data[1054] <= 14'h0429;
  filter_in_data[1055] <= 14'h0439;
  filter_in_data[1056] <= 14'h0449;
  filter_in_data[1057] <= 14'h0459;
  filter_in_data[1058] <= 14'h0469;
  filter_in_data[1059] <= 14'h0479;
  filter_in_data[1060] <= 14'h0489;
  filter_in_data[1061] <= 14'h0499;
  filter_in_data[1062] <= 14'h04a9;
  filter_in_data[1063] <= 14'h04b9;
  filter_in_data[1064] <= 14'h04c9;
  filter_in_data[1065] <= 14'h04d9;
  filter_in_data[1066] <= 14'h04e9;
  filter_in_data[1067] <= 14'h04f9;
  filter_in_data[1068] <= 14'h0509;
  filter_in_data[1069] <= 14'h0519;
  filter_in_data[1070] <= 14'h0529;
  filter_in_data[1071] <= 14'h0539;
  filter_in_data[1072] <= 14'h0549;
  filter_in_data[1073] <= 14'h0559;
  filter_in_data[1074] <= 14'h0569;
  filter_in_data[1075] <= 14'h0579;
  filter_in_data[1076] <= 14'h0589;
  filter_in_data[1077] <= 14'h0599;
  filter_in_data[1078] <= 14'h05a9;
  filter_in_data[1079] <= 14'h05b9;
  filter_in_data[1080] <= 14'h05c9;
  filter_in_data[1081] <= 14'h05d9;
  filter_in_data[1082] <= 14'h05e9;
  filter_in_data[1083] <= 14'h05f9;
  filter_in_data[1084] <= 14'h060a;
  filter_in_data[1085] <= 14'h061a;
  filter_in_data[1086] <= 14'h062a;
  filter_in_data[1087] <= 14'h063a;
  filter_in_data[1088] <= 14'h064a;
  filter_in_data[1089] <= 14'h065a;
  filter_in_data[1090] <= 14'h066a;
  filter_in_data[1091] <= 14'h067a;
  filter_in_data[1092] <= 14'h068a;
  filter_in_data[1093] <= 14'h069a;
  filter_in_data[1094] <= 14'h06aa;
  filter_in_data[1095] <= 14'h06ba;
  filter_in_data[1096] <= 14'h06ca;
  filter_in_data[1097] <= 14'h06da;
  filter_in_data[1098] <= 14'h06ea;
  filter_in_data[1099] <= 14'h06fa;
  filter_in_data[1100] <= 14'h070a;
  filter_in_data[1101] <= 14'h071a;
  filter_in_data[1102] <= 14'h072a;
  filter_in_data[1103] <= 14'h073a;
  filter_in_data[1104] <= 14'h074a;
  filter_in_data[1105] <= 14'h075a;
  filter_in_data[1106] <= 14'h076a;
  filter_in_data[1107] <= 14'h077a;
  filter_in_data[1108] <= 14'h078a;
  filter_in_data[1109] <= 14'h079a;
  filter_in_data[1110] <= 14'h07aa;
  filter_in_data[1111] <= 14'h07ba;
  filter_in_data[1112] <= 14'h07ca;
  filter_in_data[1113] <= 14'h07da;
  filter_in_data[1114] <= 14'h07ea;
  filter_in_data[1115] <= 14'h07fa;
  filter_in_data[1116] <= 14'h080a;
  filter_in_data[1117] <= 14'h081a;
  filter_in_data[1118] <= 14'h082a;
  filter_in_data[1119] <= 14'h083a;
  filter_in_data[1120] <= 14'h084a;
  filter_in_data[1121] <= 14'h085a;
  filter_in_data[1122] <= 14'h086a;
  filter_in_data[1123] <= 14'h087a;
  filter_in_data[1124] <= 14'h088a;
  filter_in_data[1125] <= 14'h089a;
  filter_in_data[1126] <= 14'h08aa;
  filter_in_data[1127] <= 14'h08ba;
  filter_in_data[1128] <= 14'h08ca;
  filter_in_data[1129] <= 14'h08da;
  filter_in_data[1130] <= 14'h08ea;
  filter_in_data[1131] <= 14'h08fa;
  filter_in_data[1132] <= 14'h090a;
  filter_in_data[1133] <= 14'h091a;
  filter_in_data[1134] <= 14'h092a;
  filter_in_data[1135] <= 14'h093a;
  filter_in_data[1136] <= 14'h094a;
  filter_in_data[1137] <= 14'h095a;
  filter_in_data[1138] <= 14'h096a;
  filter_in_data[1139] <= 14'h097a;
  filter_in_data[1140] <= 14'h098a;
  filter_in_data[1141] <= 14'h099a;
  filter_in_data[1142] <= 14'h09aa;
  filter_in_data[1143] <= 14'h09ba;
  filter_in_data[1144] <= 14'h09ca;
  filter_in_data[1145] <= 14'h09da;
  filter_in_data[1146] <= 14'h09ea;
  filter_in_data[1147] <= 14'h09fa;
  filter_in_data[1148] <= 14'h0a0b;
  filter_in_data[1149] <= 14'h0a1b;
  filter_in_data[1150] <= 14'h0a2b;
  filter_in_data[1151] <= 14'h0a3b;
  filter_in_data[1152] <= 14'h0a4b;
  filter_in_data[1153] <= 14'h0a5b;
  filter_in_data[1154] <= 14'h0a6b;
  filter_in_data[1155] <= 14'h0a7b;
  filter_in_data[1156] <= 14'h0a8b;
  filter_in_data[1157] <= 14'h0a9b;
  filter_in_data[1158] <= 14'h0aab;
  filter_in_data[1159] <= 14'h0abb;
  filter_in_data[1160] <= 14'h0acb;
  filter_in_data[1161] <= 14'h0adb;
  filter_in_data[1162] <= 14'h0aeb;
  filter_in_data[1163] <= 14'h0afb;
  filter_in_data[1164] <= 14'h0b0b;
  filter_in_data[1165] <= 14'h0b1b;
  filter_in_data[1166] <= 14'h0b2b;
  filter_in_data[1167] <= 14'h0b3b;
  filter_in_data[1168] <= 14'h0b4b;
  filter_in_data[1169] <= 14'h0b5b;
  filter_in_data[1170] <= 14'h0b6b;
  filter_in_data[1171] <= 14'h0b7b;
  filter_in_data[1172] <= 14'h0b8b;
  filter_in_data[1173] <= 14'h0b9b;
  filter_in_data[1174] <= 14'h0bab;
  filter_in_data[1175] <= 14'h0bbb;
  filter_in_data[1176] <= 14'h0bcb;
  filter_in_data[1177] <= 14'h0bdb;
  filter_in_data[1178] <= 14'h0beb;
  filter_in_data[1179] <= 14'h0bfb;
  filter_in_data[1180] <= 14'h0c0b;
  filter_in_data[1181] <= 14'h0c1b;
  filter_in_data[1182] <= 14'h0c2b;
  filter_in_data[1183] <= 14'h0c3b;
  filter_in_data[1184] <= 14'h0c4b;
  filter_in_data[1185] <= 14'h0c5b;
  filter_in_data[1186] <= 14'h0c6b;
  filter_in_data[1187] <= 14'h0c7b;
  filter_in_data[1188] <= 14'h0c8b;
  filter_in_data[1189] <= 14'h0c9b;
  filter_in_data[1190] <= 14'h0cab;
  filter_in_data[1191] <= 14'h0cbb;
  filter_in_data[1192] <= 14'h0ccb;
  filter_in_data[1193] <= 14'h0cdb;
  filter_in_data[1194] <= 14'h0ceb;
  filter_in_data[1195] <= 14'h0cfb;
  filter_in_data[1196] <= 14'h0d0b;
  filter_in_data[1197] <= 14'h0d1b;
  filter_in_data[1198] <= 14'h0d2b;
  filter_in_data[1199] <= 14'h0d3b;
  filter_in_data[1200] <= 14'h0d4b;
  filter_in_data[1201] <= 14'h0d5b;
  filter_in_data[1202] <= 14'h0d6b;
  filter_in_data[1203] <= 14'h0d7b;
  filter_in_data[1204] <= 14'h0d8b;
  filter_in_data[1205] <= 14'h0d9b;
  filter_in_data[1206] <= 14'h0dab;
  filter_in_data[1207] <= 14'h0dbb;
  filter_in_data[1208] <= 14'h0dcb;
  filter_in_data[1209] <= 14'h0ddb;
  filter_in_data[1210] <= 14'h0deb;
  filter_in_data[1211] <= 14'h0dfb;
  filter_in_data[1212] <= 14'h0e0c;
  filter_in_data[1213] <= 14'h0e1c;
  filter_in_data[1214] <= 14'h0e2c;
  filter_in_data[1215] <= 14'h0e3c;
  filter_in_data[1216] <= 14'h0e4c;
  filter_in_data[1217] <= 14'h0e5c;
  filter_in_data[1218] <= 14'h0e6c;
  filter_in_data[1219] <= 14'h0e7c;
  filter_in_data[1220] <= 14'h0e8c;
  filter_in_data[1221] <= 14'h0e9c;
  filter_in_data[1222] <= 14'h0eac;
  filter_in_data[1223] <= 14'h0ebc;
  filter_in_data[1224] <= 14'h0ecc;
  filter_in_data[1225] <= 14'h0edc;
  filter_in_data[1226] <= 14'h0eec;
  filter_in_data[1227] <= 14'h0efc;
  filter_in_data[1228] <= 14'h0f0c;
  filter_in_data[1229] <= 14'h0f1c;
  filter_in_data[1230] <= 14'h0f2c;
  filter_in_data[1231] <= 14'h0f3c;
  filter_in_data[1232] <= 14'h0f4c;
  filter_in_data[1233] <= 14'h0f5c;
  filter_in_data[1234] <= 14'h0f6c;
  filter_in_data[1235] <= 14'h0f7c;
  filter_in_data[1236] <= 14'h0f8c;
  filter_in_data[1237] <= 14'h0f9c;
  filter_in_data[1238] <= 14'h0fac;
  filter_in_data[1239] <= 14'h0fbc;
  filter_in_data[1240] <= 14'h0fcc;
  filter_in_data[1241] <= 14'h0fdc;
  filter_in_data[1242] <= 14'h0fec;
  filter_in_data[1243] <= 14'h0ffc;
  filter_in_data[1244] <= 14'h100c;
  filter_in_data[1245] <= 14'h101c;
  filter_in_data[1246] <= 14'h102c;
  filter_in_data[1247] <= 14'h103c;
  filter_in_data[1248] <= 14'h104c;
  filter_in_data[1249] <= 14'h105c;
  filter_in_data[1250] <= 14'h106c;
  filter_in_data[1251] <= 14'h107c;
  filter_in_data[1252] <= 14'h108c;
  filter_in_data[1253] <= 14'h109c;
  filter_in_data[1254] <= 14'h10ac;
  filter_in_data[1255] <= 14'h10bc;
  filter_in_data[1256] <= 14'h10cc;
  filter_in_data[1257] <= 14'h10dc;
  filter_in_data[1258] <= 14'h10ec;
  filter_in_data[1259] <= 14'h10fc;
  filter_in_data[1260] <= 14'h110c;
  filter_in_data[1261] <= 14'h111c;
  filter_in_data[1262] <= 14'h112c;
  filter_in_data[1263] <= 14'h113c;
  filter_in_data[1264] <= 14'h114c;
  filter_in_data[1265] <= 14'h115c;
  filter_in_data[1266] <= 14'h116c;
  filter_in_data[1267] <= 14'h117c;
  filter_in_data[1268] <= 14'h118c;
  filter_in_data[1269] <= 14'h119c;
  filter_in_data[1270] <= 14'h11ac;
  filter_in_data[1271] <= 14'h11bc;
  filter_in_data[1272] <= 14'h11cc;
  filter_in_data[1273] <= 14'h11dc;
  filter_in_data[1274] <= 14'h11ec;
  filter_in_data[1275] <= 14'h11fc;
  filter_in_data[1276] <= 14'h120d;
  filter_in_data[1277] <= 14'h121d;
  filter_in_data[1278] <= 14'h122d;
  filter_in_data[1279] <= 14'h123d;
  filter_in_data[1280] <= 14'h124d;
  filter_in_data[1281] <= 14'h125d;
  filter_in_data[1282] <= 14'h126d;
  filter_in_data[1283] <= 14'h127d;
  filter_in_data[1284] <= 14'h128d;
  filter_in_data[1285] <= 14'h129d;
  filter_in_data[1286] <= 14'h12ad;
  filter_in_data[1287] <= 14'h12bd;
  filter_in_data[1288] <= 14'h12cd;
  filter_in_data[1289] <= 14'h12dd;
  filter_in_data[1290] <= 14'h12ed;
  filter_in_data[1291] <= 14'h12fd;
  filter_in_data[1292] <= 14'h130d;
  filter_in_data[1293] <= 14'h131d;
  filter_in_data[1294] <= 14'h132d;
  filter_in_data[1295] <= 14'h133d;
  filter_in_data[1296] <= 14'h134d;
  filter_in_data[1297] <= 14'h135d;
  filter_in_data[1298] <= 14'h136d;
  filter_in_data[1299] <= 14'h137d;
  filter_in_data[1300] <= 14'h138d;
  filter_in_data[1301] <= 14'h139d;
  filter_in_data[1302] <= 14'h13ad;
  filter_in_data[1303] <= 14'h13bd;
  filter_in_data[1304] <= 14'h13cd;
  filter_in_data[1305] <= 14'h13dd;
  filter_in_data[1306] <= 14'h13ed;
  filter_in_data[1307] <= 14'h13fd;
  filter_in_data[1308] <= 14'h140d;
  filter_in_data[1309] <= 14'h141d;
  filter_in_data[1310] <= 14'h142d;
  filter_in_data[1311] <= 14'h143d;
  filter_in_data[1312] <= 14'h144d;
  filter_in_data[1313] <= 14'h145d;
  filter_in_data[1314] <= 14'h146d;
  filter_in_data[1315] <= 14'h147d;
  filter_in_data[1316] <= 14'h148d;
  filter_in_data[1317] <= 14'h149d;
  filter_in_data[1318] <= 14'h14ad;
  filter_in_data[1319] <= 14'h14bd;
  filter_in_data[1320] <= 14'h14cd;
  filter_in_data[1321] <= 14'h14dd;
  filter_in_data[1322] <= 14'h14ed;
  filter_in_data[1323] <= 14'h14fd;
  filter_in_data[1324] <= 14'h150d;
  filter_in_data[1325] <= 14'h151d;
  filter_in_data[1326] <= 14'h152d;
  filter_in_data[1327] <= 14'h153d;
  filter_in_data[1328] <= 14'h154d;
  filter_in_data[1329] <= 14'h155d;
  filter_in_data[1330] <= 14'h156d;
  filter_in_data[1331] <= 14'h157d;
  filter_in_data[1332] <= 14'h158d;
  filter_in_data[1333] <= 14'h159d;
  filter_in_data[1334] <= 14'h15ad;
  filter_in_data[1335] <= 14'h15bd;
  filter_in_data[1336] <= 14'h15cd;
  filter_in_data[1337] <= 14'h15dd;
  filter_in_data[1338] <= 14'h15ed;
  filter_in_data[1339] <= 14'h15fd;
  filter_in_data[1340] <= 14'h160e;
  filter_in_data[1341] <= 14'h161e;
  filter_in_data[1342] <= 14'h162e;
  filter_in_data[1343] <= 14'h163e;
  filter_in_data[1344] <= 14'h164e;
  filter_in_data[1345] <= 14'h165e;
  filter_in_data[1346] <= 14'h166e;
  filter_in_data[1347] <= 14'h167e;
  filter_in_data[1348] <= 14'h168e;
  filter_in_data[1349] <= 14'h169e;
  filter_in_data[1350] <= 14'h16ae;
  filter_in_data[1351] <= 14'h16be;
  filter_in_data[1352] <= 14'h16ce;
  filter_in_data[1353] <= 14'h16de;
  filter_in_data[1354] <= 14'h16ee;
  filter_in_data[1355] <= 14'h16fe;
  filter_in_data[1356] <= 14'h170e;
  filter_in_data[1357] <= 14'h171e;
  filter_in_data[1358] <= 14'h172e;
  filter_in_data[1359] <= 14'h173e;
  filter_in_data[1360] <= 14'h174e;
  filter_in_data[1361] <= 14'h175e;
  filter_in_data[1362] <= 14'h176e;
  filter_in_data[1363] <= 14'h177e;
  filter_in_data[1364] <= 14'h178e;
  filter_in_data[1365] <= 14'h179e;
  filter_in_data[1366] <= 14'h17ae;
  filter_in_data[1367] <= 14'h17be;
  filter_in_data[1368] <= 14'h17ce;
  filter_in_data[1369] <= 14'h17de;
  filter_in_data[1370] <= 14'h17ee;
  filter_in_data[1371] <= 14'h17fe;
  filter_in_data[1372] <= 14'h180e;
  filter_in_data[1373] <= 14'h181e;
  filter_in_data[1374] <= 14'h182e;
  filter_in_data[1375] <= 14'h183e;
  filter_in_data[1376] <= 14'h184e;
  filter_in_data[1377] <= 14'h185e;
  filter_in_data[1378] <= 14'h186e;
  filter_in_data[1379] <= 14'h187e;
  filter_in_data[1380] <= 14'h188e;
  filter_in_data[1381] <= 14'h189e;
  filter_in_data[1382] <= 14'h18ae;
  filter_in_data[1383] <= 14'h18be;
  filter_in_data[1384] <= 14'h18ce;
  filter_in_data[1385] <= 14'h18de;
  filter_in_data[1386] <= 14'h18ee;
  filter_in_data[1387] <= 14'h18fe;
  filter_in_data[1388] <= 14'h190e;
  filter_in_data[1389] <= 14'h191e;
  filter_in_data[1390] <= 14'h192e;
  filter_in_data[1391] <= 14'h193e;
  filter_in_data[1392] <= 14'h194e;
  filter_in_data[1393] <= 14'h195e;
  filter_in_data[1394] <= 14'h196e;
  filter_in_data[1395] <= 14'h197e;
  filter_in_data[1396] <= 14'h198e;
  filter_in_data[1397] <= 14'h199e;
  filter_in_data[1398] <= 14'h19ae;
  filter_in_data[1399] <= 14'h19be;
  filter_in_data[1400] <= 14'h19ce;
  filter_in_data[1401] <= 14'h19de;
  filter_in_data[1402] <= 14'h19ee;
  filter_in_data[1403] <= 14'h19fe;
  filter_in_data[1404] <= 14'h1a0f;
  filter_in_data[1405] <= 14'h1a1f;
  filter_in_data[1406] <= 14'h1a2f;
  filter_in_data[1407] <= 14'h1a3f;
  filter_in_data[1408] <= 14'h1a4f;
  filter_in_data[1409] <= 14'h1a5f;
  filter_in_data[1410] <= 14'h1a6f;
  filter_in_data[1411] <= 14'h1a7f;
  filter_in_data[1412] <= 14'h1a8f;
  filter_in_data[1413] <= 14'h1a9f;
  filter_in_data[1414] <= 14'h1aaf;
  filter_in_data[1415] <= 14'h1abf;
  filter_in_data[1416] <= 14'h1acf;
  filter_in_data[1417] <= 14'h1adf;
  filter_in_data[1418] <= 14'h1aef;
  filter_in_data[1419] <= 14'h1aff;
  filter_in_data[1420] <= 14'h1b0f;
  filter_in_data[1421] <= 14'h1b1f;
  filter_in_data[1422] <= 14'h1b2f;
  filter_in_data[1423] <= 14'h1b3f;
  filter_in_data[1424] <= 14'h1b4f;
  filter_in_data[1425] <= 14'h1b5f;
  filter_in_data[1426] <= 14'h1b6f;
  filter_in_data[1427] <= 14'h1b7f;
  filter_in_data[1428] <= 14'h1b8f;
  filter_in_data[1429] <= 14'h1b9f;
  filter_in_data[1430] <= 14'h1baf;
  filter_in_data[1431] <= 14'h1bbf;
  filter_in_data[1432] <= 14'h1bcf;
  filter_in_data[1433] <= 14'h1bdf;
  filter_in_data[1434] <= 14'h1bef;
  filter_in_data[1435] <= 14'h1bff;
  filter_in_data[1436] <= 14'h1c0f;
  filter_in_data[1437] <= 14'h1c1f;
  filter_in_data[1438] <= 14'h1c2f;
  filter_in_data[1439] <= 14'h1c3f;
  filter_in_data[1440] <= 14'h1c4f;
  filter_in_data[1441] <= 14'h1c5f;
  filter_in_data[1442] <= 14'h1c6f;
  filter_in_data[1443] <= 14'h1c7f;
  filter_in_data[1444] <= 14'h1c8f;
  filter_in_data[1445] <= 14'h1c9f;
  filter_in_data[1446] <= 14'h1caf;
  filter_in_data[1447] <= 14'h1cbf;
  filter_in_data[1448] <= 14'h1ccf;
  filter_in_data[1449] <= 14'h1cdf;
  filter_in_data[1450] <= 14'h1cef;
  filter_in_data[1451] <= 14'h1cff;
  filter_in_data[1452] <= 14'h1d0f;
  filter_in_data[1453] <= 14'h1d1f;
  filter_in_data[1454] <= 14'h1d2f;
  filter_in_data[1455] <= 14'h1d3f;
  filter_in_data[1456] <= 14'h1d4f;
  filter_in_data[1457] <= 14'h1d5f;
  filter_in_data[1458] <= 14'h1d6f;
  filter_in_data[1459] <= 14'h1d7f;
  filter_in_data[1460] <= 14'h1d8f;
  filter_in_data[1461] <= 14'h1d9f;
  filter_in_data[1462] <= 14'h1daf;
  filter_in_data[1463] <= 14'h1dbf;
  filter_in_data[1464] <= 14'h1dcf;
  filter_in_data[1465] <= 14'h1ddf;
  filter_in_data[1466] <= 14'h1def;
  filter_in_data[1467] <= 14'h1dff;
  filter_in_data[1468] <= 14'h1e10;
  filter_in_data[1469] <= 14'h1e20;
  filter_in_data[1470] <= 14'h1e30;
  filter_in_data[1471] <= 14'h1e40;
  filter_in_data[1472] <= 14'h1e50;
  filter_in_data[1473] <= 14'h1e60;
  filter_in_data[1474] <= 14'h1e70;
  filter_in_data[1475] <= 14'h1e80;
  filter_in_data[1476] <= 14'h1e90;
  filter_in_data[1477] <= 14'h1ea0;
  filter_in_data[1478] <= 14'h1eb0;
  filter_in_data[1479] <= 14'h1ec0;
  filter_in_data[1480] <= 14'h1ed0;
  filter_in_data[1481] <= 14'h1ee0;
  filter_in_data[1482] <= 14'h1ef0;
  filter_in_data[1483] <= 14'h1f00;
  filter_in_data[1484] <= 14'h1f10;
  filter_in_data[1485] <= 14'h1f20;
  filter_in_data[1486] <= 14'h1f30;
  filter_in_data[1487] <= 14'h1f40;
  filter_in_data[1488] <= 14'h1f50;
  filter_in_data[1489] <= 14'h1f60;
  filter_in_data[1490] <= 14'h1f70;
  filter_in_data[1491] <= 14'h1f80;
  filter_in_data[1492] <= 14'h1f90;
  filter_in_data[1493] <= 14'h1fa0;
  filter_in_data[1494] <= 14'h1fb0;
  filter_in_data[1495] <= 14'h1fc0;
  filter_in_data[1496] <= 14'h1fd0;
  filter_in_data[1497] <= 14'h1fe0;
  filter_in_data[1498] <= 14'h1ff0;
  filter_in_data[1499] <= 14'h1fff;
  filter_in_data[1500] <= 14'h0000;
  filter_in_data[1501] <= 14'h0000;
  filter_in_data[1502] <= 14'h0000;
  filter_in_data[1503] <= 14'h0000;
  filter_in_data[1504] <= 14'h0000;
  filter_in_data[1505] <= 14'h0000;
  filter_in_data[1506] <= 14'h0000;
  filter_in_data[1507] <= 14'h0000;
  filter_in_data[1508] <= 14'h0000;
  filter_in_data[1509] <= 14'h0000;
  filter_in_data[1510] <= 14'h0000;
  filter_in_data[1511] <= 14'h0000;
  filter_in_data[1512] <= 14'h0000;
  filter_in_data[1513] <= 14'h0000;
  filter_in_data[1514] <= 14'h0000;
  filter_in_data[1515] <= 14'h0000;
  filter_in_data[1516] <= 14'h0000;
  filter_in_data[1517] <= 14'h0000;
  filter_in_data[1518] <= 14'h0000;
  filter_in_data[1519] <= 14'h0000;
  filter_in_data[1520] <= 14'h0000;
  filter_in_data[1521] <= 14'h0000;
  filter_in_data[1522] <= 14'h0000;
  filter_in_data[1523] <= 14'h0000;
  filter_in_data[1524] <= 14'h0000;
  filter_in_data[1525] <= 14'h0000;
  filter_in_data[1526] <= 14'h0000;
  filter_in_data[1527] <= 14'h0000;
  filter_in_data[1528] <= 14'h0000;
  filter_in_data[1529] <= 14'h0000;
  filter_in_data[1530] <= 14'h0000;
  filter_in_data[1531] <= 14'h0000;
  filter_in_data[1532] <= 14'h0000;
  filter_in_data[1533] <= 14'h0000;
  filter_in_data[1534] <= 14'h0000;
  filter_in_data[1535] <= 14'h0000;
  filter_in_data[1536] <= 14'h0000;
  filter_in_data[1537] <= 14'h0000;
  filter_in_data[1538] <= 14'h0000;
  filter_in_data[1539] <= 14'h0000;
  filter_in_data[1540] <= 14'h0000;
  filter_in_data[1541] <= 14'h0000;
  filter_in_data[1542] <= 14'h0000;
  filter_in_data[1543] <= 14'h0000;
  filter_in_data[1544] <= 14'h0000;
  filter_in_data[1545] <= 14'h0000;
  filter_in_data[1546] <= 14'h0000;
  filter_in_data[1547] <= 14'h0000;
  filter_in_data[1548] <= 14'h0000;
  filter_in_data[1549] <= 14'h0000;
  filter_in_data[1550] <= 14'h0000;
  filter_in_data[1551] <= 14'h0000;
  filter_in_data[1552] <= 14'h0000;
  filter_in_data[1553] <= 14'h0000;
  filter_in_data[1554] <= 14'h0000;
  filter_in_data[1555] <= 14'h0000;
  filter_in_data[1556] <= 14'h0000;
  filter_in_data[1557] <= 14'h0000;
  filter_in_data[1558] <= 14'h0000;
  filter_in_data[1559] <= 14'h0000;
  filter_in_data[1560] <= 14'h0000;
  filter_in_data[1561] <= 14'h0000;
  filter_in_data[1562] <= 14'h0000;
  filter_in_data[1563] <= 14'h0000;
  filter_in_data[1564] <= 14'h0000;
  filter_in_data[1565] <= 14'h0000;
  filter_in_data[1566] <= 14'h0000;
  filter_in_data[1567] <= 14'h0000;
  filter_in_data[1568] <= 14'h0000;
  filter_in_data[1569] <= 14'h0000;
  filter_in_data[1570] <= 14'h0000;
  filter_in_data[1571] <= 14'h0000;
  filter_in_data[1572] <= 14'h0000;
  filter_in_data[1573] <= 14'h0000;
  filter_in_data[1574] <= 14'h0000;
  filter_in_data[1575] <= 14'h0000;
  filter_in_data[1576] <= 14'h0000;
  filter_in_data[1577] <= 14'h0000;
  filter_in_data[1578] <= 14'h0000;
  filter_in_data[1579] <= 14'h0000;
  filter_in_data[1580] <= 14'h0000;
  filter_in_data[1581] <= 14'h0000;
  filter_in_data[1582] <= 14'h0000;
  filter_in_data[1583] <= 14'h0000;
  filter_in_data[1584] <= 14'h0000;
  filter_in_data[1585] <= 14'h0000;
  filter_in_data[1586] <= 14'h0000;
  filter_in_data[1587] <= 14'h0000;
  filter_in_data[1588] <= 14'h0000;
  filter_in_data[1589] <= 14'h0000;
  filter_in_data[1590] <= 14'h0000;
  filter_in_data[1591] <= 14'h0000;
  filter_in_data[1592] <= 14'h0000;
  filter_in_data[1593] <= 14'h0000;
  filter_in_data[1594] <= 14'h0000;
  filter_in_data[1595] <= 14'h0000;
  filter_in_data[1596] <= 14'h0000;
  filter_in_data[1597] <= 14'h0000;
  filter_in_data[1598] <= 14'h0000;
  filter_in_data[1599] <= 14'h0000;
  filter_in_data[1600] <= 14'h0000;
  filter_in_data[1601] <= 14'h0000;
  filter_in_data[1602] <= 14'h0000;
  filter_in_data[1603] <= 14'h0000;
  filter_in_data[1604] <= 14'h0000;
  filter_in_data[1605] <= 14'h0000;
  filter_in_data[1606] <= 14'h0000;
  filter_in_data[1607] <= 14'h0000;
  filter_in_data[1608] <= 14'h0000;
  filter_in_data[1609] <= 14'h0000;
  filter_in_data[1610] <= 14'h0000;
  filter_in_data[1611] <= 14'h0000;
  filter_in_data[1612] <= 14'h0000;
  filter_in_data[1613] <= 14'h0000;
  filter_in_data[1614] <= 14'h0000;
  filter_in_data[1615] <= 14'h0000;
  filter_in_data[1616] <= 14'h0000;
  filter_in_data[1617] <= 14'h0000;
  filter_in_data[1618] <= 14'h0000;
  filter_in_data[1619] <= 14'h1fff;
  filter_in_data[1620] <= 14'h1fff;
  filter_in_data[1621] <= 14'h1fff;
  filter_in_data[1622] <= 14'h1fff;
  filter_in_data[1623] <= 14'h1ffe;
  filter_in_data[1624] <= 14'h1ffa;
  filter_in_data[1625] <= 14'h1ff4;
  filter_in_data[1626] <= 14'h1fea;
  filter_in_data[1627] <= 14'h1fda;
  filter_in_data[1628] <= 14'h1fc3;
  filter_in_data[1629] <= 14'h1fa3;
  filter_in_data[1630] <= 14'h1f79;
  filter_in_data[1631] <= 14'h1f40;
  filter_in_data[1632] <= 14'h1ef9;
  filter_in_data[1633] <= 14'h1e9e;
  filter_in_data[1634] <= 14'h1e2f;
  filter_in_data[1635] <= 14'h1da8;
  filter_in_data[1636] <= 14'h1d05;
  filter_in_data[1637] <= 14'h1c46;
  filter_in_data[1638] <= 14'h1b65;
  filter_in_data[1639] <= 14'h1a60;
  filter_in_data[1640] <= 14'h1935;
  filter_in_data[1641] <= 14'h17e2;
  filter_in_data[1642] <= 14'h1663;
  filter_in_data[1643] <= 14'h14b7;
  filter_in_data[1644] <= 14'h12dc;
  filter_in_data[1645] <= 14'h10d3;
  filter_in_data[1646] <= 14'h0e9a;
  filter_in_data[1647] <= 14'h0c33;
  filter_in_data[1648] <= 14'h099e;
  filter_in_data[1649] <= 14'h06e0;
  filter_in_data[1650] <= 14'h03fb;
  filter_in_data[1651] <= 14'h00f5;
  filter_in_data[1652] <= 14'h3dd4;
  filter_in_data[1653] <= 14'h3aa0;
  filter_in_data[1654] <= 14'h3763;
  filter_in_data[1655] <= 14'h3426;
  filter_in_data[1656] <= 14'h30f6;
  filter_in_data[1657] <= 14'h2de0;
  filter_in_data[1658] <= 14'h2af3;
  filter_in_data[1659] <= 14'h283d;
  filter_in_data[1660] <= 14'h25cf;
  filter_in_data[1661] <= 14'h23b9;
  filter_in_data[1662] <= 14'h220b;
  filter_in_data[1663] <= 14'h20d5;
  filter_in_data[1664] <= 14'h2024;
  filter_in_data[1665] <= 14'h2007;
  filter_in_data[1666] <= 14'h2088;
  filter_in_data[1667] <= 14'h21ae;
  filter_in_data[1668] <= 14'h237d;
  filter_in_data[1669] <= 14'h25f6;
  filter_in_data[1670] <= 14'h2914;
  filter_in_data[1671] <= 14'h2ccd;
  filter_in_data[1672] <= 14'h3111;
  filter_in_data[1673] <= 14'h35cc;
  filter_in_data[1674] <= 14'h3ae3;
  filter_in_data[1675] <= 14'h0036;
  filter_in_data[1676] <= 14'h059f;
  filter_in_data[1677] <= 14'h0af6;
  filter_in_data[1678] <= 14'h100f;
  filter_in_data[1679] <= 14'h14bb;
  filter_in_data[1680] <= 14'h18ce;
  filter_in_data[1681] <= 14'h1c1a;
  filter_in_data[1682] <= 14'h1e78;
  filter_in_data[1683] <= 14'h1fc5;
  filter_in_data[1684] <= 14'h1fe9;
  filter_in_data[1685] <= 14'h1ed4;
  filter_in_data[1686] <= 14'h1c81;
  filter_in_data[1687] <= 14'h18fc;
  filter_in_data[1688] <= 14'h145d;
  filter_in_data[1689] <= 14'h0ecb;
  filter_in_data[1690] <= 14'h087d;
  filter_in_data[1691] <= 14'h01b4;
  filter_in_data[1692] <= 14'h3abf;
  filter_in_data[1693] <= 14'h33f3;
  filter_in_data[1694] <= 14'h2da9;
  filter_in_data[1695] <= 14'h2839;
  filter_in_data[1696] <= 14'h23f7;
  filter_in_data[1697] <= 14'h2128;
  filter_in_data[1698] <= 14'h2005;
  filter_in_data[1699] <= 14'h20ad;
  filter_in_data[1700] <= 14'h2329;
  filter_in_data[1701] <= 14'h2763;
  filter_in_data[1702] <= 14'h2d2b;
  filter_in_data[1703] <= 14'h3431;
  filter_in_data[1704] <= 14'h3c0e;
  filter_in_data[1705] <= 14'h0444;
  filter_in_data[1706] <= 14'h0c49;
  filter_in_data[1707] <= 14'h138e;
  filter_in_data[1708] <= 14'h1988;
  filter_in_data[1709] <= 14'h1dbf;
  filter_in_data[1710] <= 14'h1fd3;
  filter_in_data[1711] <= 14'h1f8a;
  filter_in_data[1712] <= 14'h1cd6;
  filter_in_data[1713] <= 14'h17da;
  filter_in_data[1714] <= 14'h10e8;
  filter_in_data[1715] <= 14'h0883;
  filter_in_data[1716] <= 14'h3f52;
  filter_in_data[1717] <= 14'h3619;
  filter_in_data[1718] <= 14'h2da4;
  filter_in_data[1719] <= 14'h26ba;
  filter_in_data[1720] <= 14'h2207;
  filter_in_data[1721] <= 14'h200b;
  filter_in_data[1722] <= 14'h210b;
  filter_in_data[1723] <= 14'h2505;
  filter_in_data[1724] <= 14'h2baa;
  filter_in_data[1725] <= 14'h3465;
  filter_in_data[1726] <= 14'h3e61;
  filter_in_data[1727] <= 14'h08a0;
  filter_in_data[1728] <= 14'h120e;
  filter_in_data[1729] <= 14'h19a2;
  filter_in_data[1730] <= 14'h1e7b;
  filter_in_data[1731] <= 14'h1ffd;
  filter_in_data[1732] <= 14'h1de5;
  filter_in_data[1733] <= 14'h1857;
  filter_in_data[1734] <= 14'h0fe5;
  filter_in_data[1735] <= 14'h057b;
  filter_in_data[1736] <= 14'h3a52;
  filter_in_data[1737] <= 14'h2fc4;
  filter_in_data[1738] <= 14'h2729;
  filter_in_data[1739] <= 14'h21a6;
  filter_in_data[1740] <= 14'h2007;
  filter_in_data[1741] <= 14'h2299;
  filter_in_data[1742] <= 14'h2921;
  filter_in_data[1743] <= 14'h32d1;
  filter_in_data[1744] <= 14'h3e67;
  filter_in_data[1745] <= 14'h0a4d;
  filter_in_data[1746] <= 14'h14d3;
  filter_in_data[1747] <= 14'h1c68;
  filter_in_data[1748] <= 14'h1fdd;
  filter_in_data[1749] <= 14'h1e97;
  filter_in_data[1750] <= 14'h18ab;
  filter_in_data[1751] <= 14'h0ee7;
  filter_in_data[1752] <= 14'h02bd;
  filter_in_data[1753] <= 14'h360d;
  filter_in_data[1754] <= 14'h2ae1;
  filter_in_data[1755] <= 14'h2314;
  filter_in_data[1756] <= 14'h2004;
  filter_in_data[1757] <= 14'h2250;
  filter_in_data[1758] <= 14'h29b1;
  filter_in_data[1759] <= 14'h34fa;
  filter_in_data[1760] <= 14'h0247;
  filter_in_data[1761] <= 14'h0f42;
  filter_in_data[1762] <= 14'h1993;
  filter_in_data[1763] <= 14'h1f47;
  filter_in_data[1764] <= 14'h1f37;
  filter_in_data[1765] <= 14'h1949;
  filter_in_data[1766] <= 14'h0e7f;
  filter_in_data[1767] <= 14'h00d7;
  filter_in_data[1768] <= 14'h32ee;
  filter_in_data[1769] <= 14'h2787;
  filter_in_data[1770] <= 14'h20f9;
  filter_in_data[1771] <= 14'h20b2;
  filter_in_data[1772] <= 14'h26df;
  filter_in_data[1773] <= 14'h3256;
  filter_in_data[1774] <= 14'h00c3;
  filter_in_data[1775] <= 14'h0f1c;
  filter_in_data[1776] <= 14'h1a44;
  filter_in_data[1777] <= 14'h1fb7;
  filter_in_data[1778] <= 14'h1e23;
  filter_in_data[1779] <= 14'h15c3;
  filter_in_data[1780] <= 14'h0860;
  filter_in_data[1781] <= 14'h38fa;
  filter_in_data[1782] <= 14'h2b22;
  filter_in_data[1783] <= 14'h2226;
  filter_in_data[1784] <= 14'h2042;
  filter_in_data[1785] <= 14'h260b;
  filter_in_data[1786] <= 14'h323a;
  filter_in_data[1787] <= 14'h01e4;
  filter_in_data[1788] <= 14'h112b;
  filter_in_data[1789] <= 14'h1c2b;
  filter_in_data[1790] <= 14'h1fff;
  filter_in_data[1791] <= 14'h1b88;
  filter_in_data[1792] <= 14'h0fd0;
  filter_in_data[1793] <= 14'h3fd4;
  filter_in_data[1794] <= 14'h2fcf;
  filter_in_data[1795] <= 14'h241b;
  filter_in_data[1796] <= 14'h2001;
  filter_in_data[1797] <= 14'h24c6;
  filter_in_data[1798] <= 14'h3137;
  filter_in_data[1799] <= 14'h01ea;
  filter_in_data[1800] <= 14'h1227;
  filter_in_data[1801] <= 14'h1d33;
  filter_in_data[1802] <= 14'h1fbd;
  filter_in_data[1803] <= 14'h18e2;
  filter_in_data[1804] <= 14'h0a89;
  filter_in_data[1805] <= 14'h38ee;
  filter_in_data[1806] <= 14'h2967;
  filter_in_data[1807] <= 14'h20ca;
  filter_in_data[1808] <= 14'h21e2;
  filter_in_data[1809] <= 14'h2c7e;
  filter_in_data[1810] <= 14'h3d5e;
  filter_in_data[1811] <= 14'h0f2c;
  filter_in_data[1812] <= 14'h1c1f;
  filter_in_data[1813] <= 14'h1fe3;
  filter_in_data[1814] <= 14'h1914;
  filter_in_data[1815] <= 14'h09d4;
  filter_in_data[1816] <= 14'h372f;
  filter_in_data[1817] <= 14'h2778;
  filter_in_data[1818] <= 14'h2029;
  filter_in_data[1819] <= 14'h23ed;
  filter_in_data[1820] <= 14'h3199;
  filter_in_data[1821] <= 14'h0474;
  filter_in_data[1822] <= 14'h15ca;
  filter_in_data[1823] <= 14'h1f4d;
  filter_in_data[1824] <= 14'h1d66;
  filter_in_data[1825] <= 14'h109f;
  filter_in_data[1826] <= 14'h3d98;
  filter_in_data[1827] <= 14'h2b64;
  filter_in_data[1828] <= 14'h20f2;
  filter_in_data[1829] <= 14'h225e;
  filter_in_data[1830] <= 14'h2f44;
  filter_in_data[1831] <= 14'h02c1;
  filter_in_data[1832] <= 14'h153d;
  filter_in_data[1833] <= 14'h1f59;
  filter_in_data[1834] <= 14'h1ce9;
  filter_in_data[1835] <= 14'h0ec1;
  filter_in_data[1836] <= 14'h3a83;
  filter_in_data[1837] <= 14'h2874;
  filter_in_data[1838] <= 14'h201f;
  filter_in_data[1839] <= 14'h2522;
  filter_in_data[1840] <= 14'h358b;
  filter_in_data[1841] <= 14'h0a7b;
  filter_in_data[1842] <= 14'h1afc;
  filter_in_data[1843] <= 14'h1fd3;
  filter_in_data[1844] <= 14'h16bb;
  filter_in_data[1845] <= 14'h038e;
  filter_in_data[1846] <= 14'h2eb9;
  filter_in_data[1847] <= 14'h2195;
  filter_in_data[1848] <= 14'h2230;
  filter_in_data[1849] <= 14'h306d;
  filter_in_data[1850] <= 14'h05e7;
  filter_in_data[1851] <= 14'h18b5;
  filter_in_data[1852] <= 14'h1fff;
  filter_in_data[1853] <= 14'h1830;
  filter_in_data[1854] <= 14'h04d2;
  filter_in_data[1855] <= 14'h2f12;
  filter_in_data[1856] <= 14'h2172;
  filter_in_data[1857] <= 14'h22b2;
  filter_in_data[1858] <= 14'h3260;
  filter_in_data[1859] <= 14'h08e0;
  filter_in_data[1860] <= 14'h1b02;
  filter_in_data[1861] <= 14'h1f96;
  filter_in_data[1862] <= 14'h1420;
  filter_in_data[1863] <= 14'h3e51;
  filter_in_data[1864] <= 14'h294e;
  filter_in_data[1865] <= 14'h2008;
  filter_in_data[1866] <= 14'h277e;
  filter_in_data[1867] <= 14'h3bee;
  filter_in_data[1868] <= 14'h129a;
  filter_in_data[1869] <= 14'h1f5d;
  filter_in_data[1870] <= 14'h1b36;
  filter_in_data[1871] <= 14'h0837;
  filter_in_data[1872] <= 14'h30a6;
  filter_in_data[1873] <= 14'h2180;
  filter_in_data[1874] <= 14'h234e;
  filter_in_data[1875] <= 14'h3539;
  filter_in_data[1876] <= 14'h0d4b;
  filter_in_data[1877] <= 14'h1ddd;
  filter_in_data[1878] <= 14'h1d57;
  filter_in_data[1879] <= 14'h0bd9;
  filter_in_data[1880] <= 14'h3366;
  filter_in_data[1881] <= 14'h2246;
  filter_in_data[1882] <= 14'h22aa;
  filter_in_data[1883] <= 14'h3486;
  filter_in_data[1884] <= 14'h0d51;
  filter_in_data[1885] <= 14'h1e24;
  filter_in_data[1886] <= 14'h1cae;
  filter_in_data[1887] <= 14'h09a6;
  filter_in_data[1888] <= 14'h309c;
  filter_in_data[1889] <= 14'h210f;
  filter_in_data[1890] <= 14'h24d2;
  filter_in_data[1891] <= 14'h39b8;
  filter_in_data[1892] <= 14'h12a9;
  filter_in_data[1893] <= 14'h1fc0;
  filter_in_data[1894] <= 14'h1875;
  filter_in_data[1895] <= 14'h014d;
  filter_in_data[1896] <= 14'h293d;
  filter_in_data[1897] <= 14'h200d;
  filter_in_data[1898] <= 14'h2bf5;
  filter_in_data[1899] <= 14'h053c;
  filter_in_data[1900] <= 14'h1b13;
  filter_in_data[1901] <= 14'h1eb6;
  filter_in_data[1902] <= 14'h0d82;
  filter_in_data[1903] <= 14'h3307;
  filter_in_data[1904] <= 14'h2167;
  filter_in_data[1905] <= 14'h24ec;
  filter_in_data[1906] <= 14'h3b55;
  filter_in_data[1907] <= 14'h1512;
  filter_in_data[1908] <= 14'h1fff;
  filter_in_data[1909] <= 14'h1434;
  filter_in_data[1910] <= 14'h39ed;
  filter_in_data[1911] <= 14'h23f5;
  filter_in_data[1912] <= 14'h2242;
  filter_in_data[1913] <= 14'h363f;
  filter_in_data[1914] <= 14'h1172;
  filter_in_data[1915] <= 14'h1fd3;
  filter_in_data[1916] <= 14'h1695;
  filter_in_data[1917] <= 14'h3c6d;
  filter_in_data[1918] <= 14'h24e5;
  filter_in_data[1919] <= 14'h21d7;
  filter_in_data[1920] <= 14'h35c4;
  filter_in_data[1921] <= 14'h1196;
  filter_in_data[1922] <= 14'h1fe7;
  filter_in_data[1923] <= 14'h157b;
  filter_in_data[1924] <= 14'h3a42;
  filter_in_data[1925] <= 14'h237c;
  filter_in_data[1926] <= 14'h2335;
  filter_in_data[1927] <= 14'h39d6;
  filter_in_data[1928] <= 14'h1573;
  filter_in_data[1929] <= 14'h1fdb;
  filter_in_data[1930] <= 14'h107c;
  filter_in_data[1931] <= 14'h33a6;
  filter_in_data[1932] <= 14'h20df;
  filter_in_data[1933] <= 14'h27b9;
  filter_in_data[1934] <= 14'h02b9;
  filter_in_data[1935] <= 14'h1b83;
  filter_in_data[1936] <= 14'h1d44;
  filter_in_data[1937] <= 14'h0652;
  filter_in_data[1938] <= 14'h29f6;
  filter_in_data[1939] <= 14'h205d;
  filter_in_data[1940] <= 14'h31ea;
  filter_in_data[1941] <= 14'h0fac;
  filter_in_data[1942] <= 14'h1fe0;
  filter_in_data[1943] <= 14'h1443;
  filter_in_data[1944] <= 14'h36d2;
  filter_in_data[1945] <= 14'h216e;
  filter_in_data[1946] <= 14'h272a;
  filter_in_data[1947] <= 14'h031b;
  filter_in_data[1948] <= 14'h1c50;
  filter_in_data[1949] <= 14'h1bfb;
  filter_in_data[1950] <= 14'h0238;
  filter_in_data[1951] <= 14'h2662;
  filter_in_data[1952] <= 14'h2208;
  filter_in_data[1953] <= 14'h395c;
  filter_in_data[1954] <= 14'h16e7;
  filter_in_data[1955] <= 14'h1f1c;
  filter_in_data[1956] <= 14'h0a1d;
  filter_in_data[1957] <= 14'h2b87;
  filter_in_data[1958] <= 14'h2053;
  filter_in_data[1959] <= 14'h3356;
  filter_in_data[1960] <= 14'h1289;
  filter_in_data[1961] <= 14'h1fe9;
  filter_in_data[1962] <= 14'h0e5b;
  filter_in_data[1963] <= 14'h2ec5;
  filter_in_data[1964] <= 14'h2005;
  filter_in_data[1965] <= 14'h30c2;
  filter_in_data[1966] <= 14'h10a0;
  filter_in_data[1967] <= 14'h1ffe;
  filter_in_data[1968] <= 14'h0f5c;
  filter_in_data[1969] <= 14'h2f3e;
  filter_in_data[1970] <= 14'h2005;
  filter_in_data[1971] <= 14'h314a;
  filter_in_data[1972] <= 14'h119f;
  filter_in_data[1973] <= 14'h1fe8;
  filter_in_data[1974] <= 14'h0d45;
  filter_in_data[1975] <= 14'h2cd5;
  filter_in_data[1976] <= 14'h2055;
  filter_in_data[1977] <= 14'h3503;
  filter_in_data[1978] <= 14'h154d;
  filter_in_data[1979] <= 14'h1f16;
  filter_in_data[1980] <= 14'h07ce;
  filter_in_data[1981] <= 14'h2823;
  filter_in_data[1982] <= 14'h2212;
  filter_in_data[1983] <= 14'h3c54;
  filter_in_data[1984] <= 14'h1a9c;
  filter_in_data[1985] <= 14'h1be9;
  filter_in_data[1986] <= 14'h3e9d;
  filter_in_data[1987] <= 14'h22cd;
  filter_in_data[1988] <= 14'h2745;
  filter_in_data[1989] <= 14'h0742;
  filter_in_data[1990] <= 14'h1f2e;
  filter_in_data[1991] <= 14'h141d;
  filter_in_data[1992] <= 14'h3255;
  filter_in_data[1993] <= 14'h2000;
  filter_in_data[1994] <= 14'h321b;
  filter_in_data[1995] <= 14'h1425;
  filter_in_data[1996] <= 14'h1f0f;
  filter_in_data[1997] <= 14'h0617;
  filter_in_data[1998] <= 14'h2604;
  filter_in_data[1999] <= 14'h2437;
  filter_in_data[2000] <= 14'h02fb;
  filter_in_data[2001] <= 14'h1e48;
  filter_in_data[2002] <= 14'h15ca;
  filter_in_data[2003] <= 14'h3363;
  filter_in_data[2004] <= 14'h2000;
  filter_in_data[2005] <= 14'h32fb;
  filter_in_data[2006] <= 14'h15ad;
  filter_in_data[2007] <= 14'h1e2c;
  filter_in_data[2008] <= 14'h01fc;
  filter_in_data[2009] <= 14'h2356;
  filter_in_data[2010] <= 14'h27d4;
  filter_in_data[2011] <= 14'h0a21;
  filter_in_data[2012] <= 14'h1fed;
  filter_in_data[2013] <= 14'h0e09;
  filter_in_data[2014] <= 14'h2a96;
  filter_in_data[2015] <= 14'h21f8;
  filter_in_data[2016] <= 14'h3f34;
  filter_in_data[2017] <= 14'h1d7b;
  filter_in_data[2018] <= 14'h164c;
  filter_in_data[2019] <= 14'h329e;
  filter_in_data[2020] <= 14'h2012;
  filter_in_data[2021] <= 14'h36a7;
  filter_in_data[2022] <= 14'h195c;
  filter_in_data[2023] <= 14'h1b24;
  filter_in_data[2024] <= 14'h397c;
  filter_in_data[2025] <= 14'h2056;
  filter_in_data[2026] <= 14'h30dc;
  filter_in_data[2027] <= 14'h156d;
  filter_in_data[2028] <= 14'h1d92;
  filter_in_data[2029] <= 14'h3e48;
  filter_in_data[2030] <= 14'h2143;
  filter_in_data[2031] <= 14'h2d90;
  filter_in_data[2032] <= 14'h12c9;
  filter_in_data[2033] <= 14'h1e90;
  filter_in_data[2034] <= 14'h00b6;
  filter_in_data[2035] <= 14'h21dc;
  filter_in_data[2036] <= 14'h2c62;
  filter_in_data[2037] <= 14'h11fa;
  filter_in_data[2038] <= 14'h1eb5;
  filter_in_data[2039] <= 14'h00bd;
  filter_in_data[2040] <= 14'h21b6;
  filter_in_data[2041] <= 14'h2d22;
  filter_in_data[2042] <= 14'h1322;
  filter_in_data[2043] <= 14'h1e1e;
  filter_in_data[2044] <= 14'h3e5b;
  filter_in_data[2045] <= 14'h20e8;
  filter_in_data[2046] <= 14'h2fef;
  filter_in_data[2047] <= 14'h160f;
  filter_in_data[2048] <= 14'h1c65;
  filter_in_data[2049] <= 14'h399b;
  filter_in_data[2050] <= 14'h2016;
  filter_in_data[2051] <= 14'h3524;
  filter_in_data[2052] <= 14'h1a21;
  filter_in_data[2053] <= 14'h18b2;
  filter_in_data[2054] <= 14'h32c6;
  filter_in_data[2055] <= 14'h2071;
  filter_in_data[2056] <= 14'h3d16;
  filter_in_data[2057] <= 14'h1e1c;
  filter_in_data[2058] <= 14'h11f9;
  filter_in_data[2059] <= 14'h2ac0;
  filter_in_data[2060] <= 14'h23a2;
  filter_in_data[2061] <= 14'h0794;
  filter_in_data[2062] <= 14'h1fff;
  filter_in_data[2063] <= 14'h077c;
  filter_in_data[2064] <= 14'h2375;
  filter_in_data[2065] <= 14'h2b68;
  filter_in_data[2066] <= 14'h133b;
  filter_in_data[2067] <= 14'h1d36;
  filter_in_data[2068] <= 14'h39a8;
  filter_in_data[2069] <= 14'h2001;
  filter_in_data[2070] <= 14'h3899;
  filter_in_data[2071] <= 14'h1ce1;
  filter_in_data[2072] <= 14'h137a;
  filter_in_data[2073] <= 14'h2b21;
  filter_in_data[2074] <= 14'h2408;
  filter_in_data[2075] <= 14'h09b0;
  filter_in_data[2076] <= 14'h1fce;
  filter_in_data[2077] <= 14'h02aa;
  filter_in_data[2078] <= 14'h2132;
  filter_in_data[2079] <= 14'h31bb;
  filter_in_data[2080] <= 14'h1988;
  filter_in_data[2081] <= 14'h1797;
  filter_in_data[2082] <= 14'h2eec;
  filter_in_data[2083] <= 14'h225e;
  filter_in_data[2084] <= 14'h06cd;
  filter_in_data[2085] <= 14'h1ff8;
  filter_in_data[2086] <= 14'h03e9;
  filter_in_data[2087] <= 14'h214e;
  filter_in_data[2088] <= 14'h322a;
  filter_in_data[2089] <= 14'h1a52;
  filter_in_data[2090] <= 14'h160a;
  filter_in_data[2091] <= 14'h2c66;
  filter_in_data[2092] <= 14'h2414;
  filter_in_data[2093] <= 14'h0b69;
  filter_in_data[2094] <= 14'h1f37;
  filter_in_data[2095] <= 14'h3d60;
  filter_in_data[2096] <= 14'h200c;
  filter_in_data[2097] <= 14'h3a02;
  filter_in_data[2098] <= 14'h1e62;
  filter_in_data[2099] <= 14'h0dd4;
  filter_in_data[2100] <= 14'h2516;
  filter_in_data[2101] <= 14'h2b8d;
  filter_in_data[2102] <= 14'h1605;
  filter_in_data[2103] <= 14'h199b;
  filter_in_data[2104] <= 14'h2fcf;
  filter_in_data[2105] <= 14'h22cb;
  filter_in_data[2106] <= 14'h09e4;
  filter_in_data[2107] <= 14'h1f4b;
  filter_in_data[2108] <= 14'h3c7d;
  filter_in_data[2109] <= 14'h2001;
  filter_in_data[2110] <= 14'h3d5e;
  filter_in_data[2111] <= 14'h1f84;
  filter_in_data[2112] <= 14'h084e;
  filter_in_data[2113] <= 14'h21eb;
  filter_in_data[2114] <= 14'h32a4;
  filter_in_data[2115] <= 14'h1bec;
  filter_in_data[2116] <= 14'h11b8;
  filter_in_data[2117] <= 14'h26ba;
  filter_in_data[2118] <= 14'h2aa3;
  filter_in_data[2119] <= 14'h1655;
  filter_in_data[2120] <= 14'h1850;
  filter_in_data[2121] <= 14'h2cba;
  filter_in_data[2122] <= 14'h255f;
  filter_in_data[2123] <= 14'h103e;
  filter_in_data[2124] <= 14'h1c63;
  filter_in_data[2125] <= 14'h32a6;
  filter_in_data[2126] <= 14'h2254;
  filter_in_data[2127] <= 14'h0aaf;
  filter_in_data[2128] <= 14'h1e92;
  filter_in_data[2129] <= 14'h37b2;
  filter_in_data[2130] <= 14'h20d4;
  filter_in_data[2131] <= 14'h0641;
  filter_in_data[2132] <= 14'h1f8c;
  filter_in_data[2133] <= 14'h3b71;
  filter_in_data[2134] <= 14'h203b;
  filter_in_data[2135] <= 14'h033b;
  filter_in_data[2136] <= 14'h1fe3;
  filter_in_data[2137] <= 14'h3db7;
  filter_in_data[2138] <= 14'h200f;
  filter_in_data[2139] <= 14'h01b8;
  filter_in_data[2140] <= 14'h1ff6;
  filter_in_data[2141] <= 14'h3e76;
  filter_in_data[2142] <= 14'h200a;
  filter_in_data[2143] <= 14'h01be;
  filter_in_data[2144] <= 14'h1ff0;
  filter_in_data[2145] <= 14'h3dab;
  filter_in_data[2146] <= 14'h201f;
  filter_in_data[2147] <= 14'h034d;
  filter_in_data[2148] <= 14'h1fc2;
  filter_in_data[2149] <= 14'h3b59;
  filter_in_data[2150] <= 14'h2078;
  filter_in_data[2151] <= 14'h065f;
  filter_in_data[2152] <= 14'h1f24;
  filter_in_data[2153] <= 14'h378f;
  filter_in_data[2154] <= 14'h217a;
  filter_in_data[2155] <= 14'h0ad7;
  filter_in_data[2156] <= 14'h1d9b;
  filter_in_data[2157] <= 14'h327a;
  filter_in_data[2158] <= 14'h23b5;
  filter_in_data[2159] <= 14'h106c;
  filter_in_data[2160] <= 14'h1a81;
  filter_in_data[2161] <= 14'h2c8a;
  filter_in_data[2162] <= 14'h27d9;
  filter_in_data[2163] <= 14'h1684;
  filter_in_data[2164] <= 14'h1529;
  filter_in_data[2165] <= 14'h268e;
  filter_in_data[2166] <= 14'h2e87;
  filter_in_data[2167] <= 14'h1c12;
  filter_in_data[2168] <= 14'h0d12;
  filter_in_data[2169] <= 14'h21cf;
  filter_in_data[2170] <= 14'h3807;
  filter_in_data[2171] <= 14'h1f94;
  filter_in_data[2172] <= 14'h0244;
  filter_in_data[2173] <= 14'h2002;
  filter_in_data[2174] <= 14'h03e6;
  filter_in_data[2175] <= 14'h1f35;
  filter_in_data[2176] <= 14'h35b8;
  filter_in_data[2177] <= 14'h22f8;
  filter_in_data[2178] <= 14'h1091;
  filter_in_data[2179] <= 14'h1956;
  filter_in_data[2180] <= 14'h29a6;
  filter_in_data[2181] <= 14'h2beb;
  filter_in_data[2182] <= 14'h1b2c;
  filter_in_data[2183] <= 14'h0d61;
  filter_in_data[2184] <= 14'h2176;
  filter_in_data[2185] <= 14'h3a85;
  filter_in_data[2186] <= 14'h1ffa;
  filter_in_data[2187] <= 14'h3cd6;
  filter_in_data[2188] <= 14'h20e9;
  filter_in_data[2189] <= 14'h0bf0;
  filter_in_data[2190] <= 14'h1ba2;
  filter_in_data[2191] <= 14'h2bf0;
  filter_in_data[2192] <= 14'h2a66;
  filter_in_data[2193] <= 14'h1aaa;
  filter_in_data[2194] <= 14'h0d45;
  filter_in_data[2195] <= 14'h2121;
  filter_in_data[2196] <= 14'h3cbc;
  filter_in_data[2197] <= 14'h1fef;
  filter_in_data[2198] <= 14'h388b;
  filter_in_data[2199] <= 14'h22a2;
  filter_in_data[2200] <= 14'h11a9;
  filter_in_data[2201] <= 14'h171c;
  filter_in_data[2202] <= 14'h260b;
  filter_in_data[2203] <= 14'h3264;
  filter_in_data[2204] <= 14'h1eff;
  filter_in_data[2205] <= 14'h01e9;
  filter_in_data[2206] <= 14'h204a;
  filter_in_data[2207] <= 14'h0a6d;
  filter_in_data[2208] <= 14'h1b93;
  filter_in_data[2209] <= 14'h2a88;
  filter_in_data[2210] <= 14'h2d2d;
  filter_in_data[2211] <= 14'h1d39;
  filter_in_data[2212] <= 14'h0696;
  filter_in_data[2213] <= 14'h2000;
  filter_in_data[2214] <= 14'h0730;
  filter_in_data[2215] <= 14'h1cd8;
  filter_in_data[2216] <= 14'h2c12;
  filter_in_data[2217] <= 14'h2c1a;
  filter_in_data[2218] <= 14'h1cf1;
  filter_in_data[2219] <= 14'h0696;
  filter_in_data[2220] <= 14'h2003;
  filter_in_data[2221] <= 14'h087e;
  filter_in_data[2222] <= 14'h1be9;
  filter_in_data[2223] <= 14'h2a09;
  filter_in_data[2224] <= 14'h2ed8;
  filter_in_data[2225] <= 14'h1e6f;
  filter_in_data[2226] <= 14'h01ea;
  filter_in_data[2227] <= 14'h209f;
  filter_in_data[2228] <= 14'h0e27;
  filter_in_data[2229] <= 14'h1806;
  filter_in_data[2230] <= 14'h2547;
  filter_in_data[2231] <= 14'h3625;
  filter_in_data[2232] <= 14'h1ff9;
  filter_in_data[2233] <= 14'h388c;
  filter_in_data[2234] <= 14'h2421;
  filter_in_data[2235] <= 14'h16d9;
  filter_in_data[2236] <= 14'h0f17;
  filter_in_data[2237] <= 14'h20a9;
  filter_in_data[2238] <= 14'h02c9;
  filter_in_data[2239] <= 14'h1db5;
  filter_in_data[2240] <= 14'h2bf1;
  filter_in_data[2241] <= 14'h2e19;
  filter_in_data[2242] <= 14'h1ea7;
  filter_in_data[2243] <= 14'h3f89;
  filter_in_data[2244] <= 14'h21a8;
  filter_in_data[2245] <= 14'h12fb;
  filter_in_data[2246] <= 14'h12a0;
  filter_in_data[2247] <= 14'h2176;
  filter_in_data[2248] <= 14'h008d;
  filter_in_data[2249] <= 14'h1e29;
  filter_in_data[2250] <= 14'h2c30;
  filter_in_data[2251] <= 14'h2ea3;
  filter_in_data[2252] <= 14'h1f14;
  filter_in_data[2253] <= 14'h3cf7;
  filter_in_data[2254] <= 14'h22f7;
  filter_in_data[2255] <= 14'h1667;
  filter_in_data[2256] <= 14'h0def;
  filter_in_data[2257] <= 14'h202b;
  filter_in_data[2258] <= 14'h07dc;
  filter_in_data[2259] <= 14'h1a60;
  filter_in_data[2260] <= 14'h25cf;
  filter_in_data[2261] <= 14'h3803;
  filter_in_data[2262] <= 14'h1fce;
  filter_in_data[2263] <= 14'h3153;
  filter_in_data[2264] <= 14'h2ac4;
  filter_in_data[2265] <= 14'h1e05;
  filter_in_data[2266] <= 14'h3f52;
  filter_in_data[2267] <= 14'h2284;
  filter_in_data[2268] <= 14'h1681;
  filter_in_data[2269] <= 14'h0caa;
  filter_in_data[2270] <= 14'h2002;
  filter_in_data[2271] <= 14'h0b92;
  filter_in_data[2272] <= 14'h1722;
  filter_in_data[2273] <= 14'h22ad;
  filter_in_data[2274] <= 14'h3f95;
  filter_in_data[2275] <= 14'h1d9c;
  filter_in_data[2276] <= 14'h292e;
  filter_in_data[2277] <= 14'h3476;
  filter_in_data[2278] <= 14'h1ff9;
  filter_in_data[2279] <= 14'h31e8;
  filter_in_data[2280] <= 14'h2b71;
  filter_in_data[2281] <= 14'h1ec6;
  filter_in_data[2282] <= 14'h3b5e;
  filter_in_data[2283] <= 14'h2515;
  filter_in_data[2284] <= 14'h1aef;
  filter_in_data[2285] <= 14'h046a;
  filter_in_data[2286] <= 14'h2166;
  filter_in_data[2287] <= 14'h1574;
  filter_in_data[2288] <= 14'h0c50;
  filter_in_data[2289] <= 14'h200a;
  filter_in_data[2290] <= 14'h0f3c;
  filter_in_data[2291] <= 14'h12b5;
  filter_in_data[2292] <= 14'h2078;
  filter_in_data[2293] <= 14'h08fe;
  filter_in_data[2294] <= 14'h178c;
  filter_in_data[2295] <= 14'h221b;
  filter_in_data[2296] <= 14'h0336;
  filter_in_data[2297] <= 14'h1af7;
  filter_in_data[2298] <= 14'h2468;
  filter_in_data[2299] <= 14'h3e2f;
  filter_in_data[2300] <= 14'h1d37;
  filter_in_data[2301] <= 14'h26ec;
  filter_in_data[2302] <= 14'h3a0d;
  filter_in_data[2303] <= 14'h1e94;
  filter_in_data[2304] <= 14'h294e;
  filter_in_data[2305] <= 14'h36d9;
  filter_in_data[2306] <= 14'h1f54;
  filter_in_data[2307] <= 14'h2b4d;
  filter_in_data[2308] <= 14'h348c;
  filter_in_data[2309] <= 14'h1fb2;
  filter_in_data[2310] <= 14'h2cc0;
  filter_in_data[2311] <= 14'h3319;
  filter_in_data[2312] <= 14'h1fd8;
  filter_in_data[2313] <= 14'h2d8c;
  filter_in_data[2314] <= 14'h3276;
  filter_in_data[2315] <= 14'h1fe2;
  filter_in_data[2316] <= 14'h2da5;
  filter_in_data[2317] <= 14'h329d;
  filter_in_data[2318] <= 14'h1fd7;
  filter_in_data[2319] <= 14'h2d0a;
  filter_in_data[2320] <= 14'h3390;
  filter_in_data[2321] <= 14'h1faf;
  filter_in_data[2322] <= 14'h2bc4;
  filter_in_data[2323] <= 14'h3555;
  filter_in_data[2324] <= 14'h1f4d;
  filter_in_data[2325] <= 14'h29e8;
  filter_in_data[2326] <= 14'h37fb;
  filter_in_data[2327] <= 14'h1e86;
  filter_in_data[2328] <= 14'h279d;
  filter_in_data[2329] <= 14'h3b8b;
  filter_in_data[2330] <= 14'h1d1e;
  filter_in_data[2331] <= 14'h251a;
  filter_in_data[2332] <= 14'h0008;
  filter_in_data[2333] <= 14'h1ad0;
  filter_in_data[2334] <= 14'h22b3;
  filter_in_data[2335] <= 14'h0560;
  filter_in_data[2336] <= 14'h1752;
  filter_in_data[2337] <= 14'h20d4;
  filter_in_data[2338] <= 14'h0b61;
  filter_in_data[2339] <= 14'h1267;
  filter_in_data[2340] <= 14'h2001;
  filter_in_data[2341] <= 14'h11af;
  filter_in_data[2342] <= 14'h0beb;
  filter_in_data[2343] <= 14'h20ce;
  filter_in_data[2344] <= 14'h17b6;
  filter_in_data[2345] <= 14'h03f2;
  filter_in_data[2346] <= 14'h23cc;
  filter_in_data[2347] <= 14'h1cac;
  filter_in_data[2348] <= 14'h3adb;
  filter_in_data[2349] <= 14'h2964;
  filter_in_data[2350] <= 14'h1f9b;
  filter_in_data[2351] <= 14'h3167;
  filter_in_data[2352] <= 14'h31b2;
  filter_in_data[2353] <= 14'h1f85;
  filter_in_data[2354] <= 14'h28c2;
  filter_in_data[2355] <= 14'h3c54;
  filter_in_data[2356] <= 14'h1b99;
  filter_in_data[2357] <= 14'h226b;
  filter_in_data[2358] <= 14'h083d;
  filter_in_data[2359] <= 14'h1382;
  filter_in_data[2360] <= 14'h2000;
  filter_in_data[2361] <= 14'h13b1;
  filter_in_data[2362] <= 14'h07bc;
  filter_in_data[2363] <= 14'h22d1;
  filter_in_data[2364] <= 14'h1c69;
  filter_in_data[2365] <= 14'h39d1;
  filter_in_data[2366] <= 14'h2b60;
  filter_in_data[2367] <= 14'h1ffe;
  filter_in_data[2368] <= 14'h2c60;
  filter_in_data[2369] <= 14'h38d7;
  filter_in_data[2370] <= 14'h1ca5;
  filter_in_data[2371] <= 14'h22c1;
  filter_in_data[2372] <= 14'h08b9;
  filter_in_data[2373] <= 14'h1203;
  filter_in_data[2374] <= 14'h202b;
  filter_in_data[2375] <= 14'h1711;
  filter_in_data[2376] <= 14'h01ea;
  filter_in_data[2377] <= 14'h2682;
  filter_in_data[2378] <= 14'h1f4c;
  filter_in_data[2379] <= 14'h3083;
  filter_in_data[2380] <= 14'h3519;
  filter_in_data[2381] <= 14'h1dcc;
  filter_in_data[2382] <= 14'h2385;
  filter_in_data[2383] <= 14'h0806;
  filter_in_data[2384] <= 14'h11bb;
  filter_in_data[2385] <= 14'h2057;
  filter_in_data[2386] <= 14'h18b3;
  filter_in_data[2387] <= 14'h3e67;
  filter_in_data[2388] <= 14'h2986;
  filter_in_data[2389] <= 14'h1ffb;
  filter_in_data[2390] <= 14'h2b0a;
  filter_in_data[2391] <= 14'h3ca2;
  filter_in_data[2392] <= 14'h1980;
  filter_in_data[2393] <= 14'h206f;
  filter_in_data[2394] <= 14'h11f0;
  filter_in_data[2395] <= 14'h06c1;
  filter_in_data[2396] <= 14'h24c7;
  filter_in_data[2397] <= 14'h1f05;
  filter_in_data[2398] <= 14'h2ffe;
  filter_in_data[2399] <= 14'h3769;
  filter_in_data[2400] <= 14'h1bfc;
  filter_in_data[2401] <= 14'h2146;
  filter_in_data[2402] <= 14'h0f5e;
  filter_in_data[2403] <= 14'h08ed;
  filter_in_data[2404] <= 14'h2408;
  filter_in_data[2405] <= 14'h1ed7;
  filter_in_data[2406] <= 14'h2fee;
  filter_in_data[2407] <= 14'h3839;
  filter_in_data[2408] <= 14'h1b2b;
  filter_in_data[2409] <= 14'h20b2;
  filter_in_data[2410] <= 14'h120e;
  filter_in_data[2411] <= 14'h051a;
  filter_in_data[2412] <= 14'h269b;
  filter_in_data[2413] <= 14'h1fd8;
  filter_in_data[2414] <= 14'h2ae1;
  filter_in_data[2415] <= 14'h3f26;
  filter_in_data[2416] <= 14'h164d;
  filter_in_data[2417] <= 14'h200e;
  filter_in_data[2418] <= 14'h18e1;
  filter_in_data[2419] <= 14'h3b0f;
  filter_in_data[2420] <= 14'h2e89;
  filter_in_data[2421] <= 14'h1ee4;
  filter_in_data[2422] <= 14'h235c;
  filter_in_data[2423] <= 14'h0c04;
  filter_in_data[2424] <= 14'h0a89;
  filter_in_data[2425] <= 14'h2432;
  filter_in_data[2426] <= 14'h1f62;
  filter_in_data[2427] <= 14'h2c4f;
  filter_in_data[2428] <= 14'h3e8c;
  filter_in_data[2429] <= 14'h15d5;
  filter_in_data[2430] <= 14'h2039;
  filter_in_data[2431] <= 14'h1abc;
  filter_in_data[2432] <= 14'h36c4;
  filter_in_data[2433] <= 14'h3385;
  filter_in_data[2434] <= 14'h1c63;
  filter_in_data[2435] <= 14'h20b0;
  filter_in_data[2436] <= 14'h1419;
  filter_in_data[2437] <= 14'h0013;
  filter_in_data[2438] <= 14'h2bdd;
  filter_in_data[2439] <= 14'h1f43;
  filter_in_data[2440] <= 14'h234a;
  filter_in_data[2441] <= 14'h0dc1;
  filter_in_data[2442] <= 14'h070c;
  filter_in_data[2443] <= 14'h273b;
  filter_in_data[2444] <= 14'h1ffd;
  filter_in_data[2445] <= 14'h262e;
  filter_in_data[2446] <= 14'h08fd;
  filter_in_data[2447] <= 14'h0b78;
  filter_in_data[2448] <= 14'h24d2;
  filter_in_data[2449] <= 14'h1fe0;
  filter_in_data[2450] <= 14'h282e;
  filter_in_data[2451] <= 14'h065f;
  filter_in_data[2452] <= 14'h0d82;
  filter_in_data[2453] <= 14'h23f2;
  filter_in_data[2454] <= 14'h1fbd;
  filter_in_data[2455] <= 14'h28b4;
  filter_in_data[2456] <= 14'h0616;
  filter_in_data[2457] <= 14'h0d55;
  filter_in_data[2458] <= 14'h2447;
  filter_in_data[2459] <= 14'h1fdd;
  filter_in_data[2460] <= 14'h279d;
  filter_in_data[2461] <= 14'h0826;
  filter_in_data[2462] <= 14'h0aee;
  filter_in_data[2463] <= 14'h25f1;
  filter_in_data[2464] <= 14'h1ffe;
  filter_in_data[2465] <= 14'h2532;
  filter_in_data[2466] <= 14'h0c6e;
  filter_in_data[2467] <= 14'h061c;
  filter_in_data[2468] <= 14'h297e;
  filter_in_data[2469] <= 14'h1f53;
  filter_in_data[2470] <= 14'h223d;
  filter_in_data[2471] <= 14'h127a;
  filter_in_data[2472] <= 14'h3ebb;
  filter_in_data[2473] <= 14'h2fbb;
  filter_in_data[2474] <= 14'h1c91;
  filter_in_data[2475] <= 14'h2028;
  filter_in_data[2476] <= 14'h1937;
  filter_in_data[2477] <= 14'h3521;
  filter_in_data[2478] <= 14'h394a;
  filter_in_data[2479] <= 14'h1630;
  filter_in_data[2480] <= 14'h2104;
  filter_in_data[2481] <= 14'h1e9b;
  filter_in_data[2482] <= 14'h2ab1;
  filter_in_data[2483] <= 14'h05ea;
  filter_in_data[2484] <= 14'h0b17;
  filter_in_data[2485] <= 14'h271e;
  filter_in_data[2486] <= 14'h1fa9;
  filter_in_data[2487] <= 14'h2256;
  filter_in_data[2488] <= 14'h1394;
  filter_in_data[2489] <= 14'h3bbd;
  filter_in_data[2490] <= 14'h33e3;
  filter_in_data[2491] <= 14'h1934;
  filter_in_data[2492] <= 14'h205a;
  filter_in_data[2493] <= 14'h1de5;
  filter_in_data[2494] <= 14'h2b7a;
  filter_in_data[2495] <= 14'h0608;
  filter_in_data[2496] <= 14'h09e3;
  filter_in_data[2497] <= 14'h28b7;
  filter_in_data[2498] <= 14'h1ef0;
  filter_in_data[2499] <= 14'h20e4;
  filter_in_data[2500] <= 14'h17e3;
  filter_in_data[2501] <= 14'h34e9;
  filter_in_data[2502] <= 14'h3bcc;
  filter_in_data[2503] <= 14'h1272;
  filter_in_data[2504] <= 14'h2392;
  filter_in_data[2505] <= 14'h1fff;
  filter_in_data[2506] <= 14'h2385;
  filter_in_data[2507] <= 14'h12c4;
  filter_in_data[2508] <= 14'h3aef;
  filter_in_data[2509] <= 14'h3660;
  filter_in_data[2510] <= 14'h1636;
  filter_in_data[2511] <= 14'h21e3;
  filter_in_data[2512] <= 14'h1fce;
  filter_in_data[2513] <= 14'h24f1;
  filter_in_data[2514] <= 14'h10f3;
  filter_in_data[2515] <= 14'h3c70;
  filter_in_data[2516] <= 14'h3592;
  filter_in_data[2517] <= 14'h1655;
  filter_in_data[2518] <= 14'h220f;
  filter_in_data[2519] <= 14'h1fea;
  filter_in_data[2520] <= 14'h23ff;
  filter_in_data[2521] <= 14'h1309;
  filter_in_data[2522] <= 14'h3947;
  filter_in_data[2523] <= 14'h394d;
  filter_in_data[2524] <= 14'h12dc;
  filter_in_data[2525] <= 14'h244b;
  filter_in_data[2526] <= 14'h1fce;
  filter_in_data[2527] <= 14'h216e;
  filter_in_data[2528] <= 14'h1853;
  filter_in_data[2529] <= 14'h31d2;
  filter_in_data[2530] <= 14'h01d8;
  filter_in_data[2531] <= 14'h0ab1;
  filter_in_data[2532] <= 14'h2a84;
  filter_in_data[2533] <= 14'h1cec;
  filter_in_data[2534] <= 14'h200b;
  filter_in_data[2535] <= 14'h1e3d;
  filter_in_data[2536] <= 14'h27e0;
  filter_in_data[2537] <= 14'h0e99;
  filter_in_data[2538] <= 14'h3cec;
  filter_in_data[2539] <= 14'h3738;
  filter_in_data[2540] <= 14'h1359;
  filter_in_data[2541] <= 14'h24c6;
  filter_in_data[2542] <= 14'h1f70;
  filter_in_data[2543] <= 14'h207c;
  filter_in_data[2544] <= 14'h1b8d;
  filter_in_data[2545] <= 14'h2bdb;
  filter_in_data[2546] <= 14'h0a4d;
  filter_in_data[2547] <= 14'h00b9;
  filter_in_data[2548] <= 14'h346f;
  filter_in_data[2549] <= 14'h14f5;
  filter_in_data[2550] <= 14'h2429;
  filter_in_data[2551] <= 14'h1f7f;
  filter_in_data[2552] <= 14'h2066;
  filter_in_data[2553] <= 14'h1c3c;
  filter_in_data[2554] <= 14'h2a26;
  filter_in_data[2555] <= 14'h0d35;
  filter_in_data[2556] <= 14'h3cbb;
  filter_in_data[2557] <= 14'h3915;
  filter_in_data[2558] <= 14'h1051;
  filter_in_data[2559] <= 14'h27fa;
  filter_in_data[2560] <= 14'h1d57;
  filter_in_data[2561] <= 14'h202b;
  filter_in_data[2562] <= 14'h1f58;
  filter_in_data[2563] <= 14'h23fe;
  filter_in_data[2564] <= 14'h1635;
  filter_in_data[2565] <= 14'h317b;
  filter_in_data[2566] <= 14'h05a9;
  filter_in_data[2567] <= 14'h0395;
  filter_in_data[2568] <= 14'h3390;
  filter_in_data[2569] <= 14'h1434;
  filter_in_data[2570] <= 14'h25b5;
  filter_in_data[2571] <= 14'h1e4a;
  filter_in_data[2572] <= 14'h200c;
  filter_in_data[2573] <= 14'h1f3d;
  filter_in_data[2574] <= 14'h23ba;
  filter_in_data[2575] <= 14'h1756;
  filter_in_data[2576] <= 14'h2f28;
  filter_in_data[2577] <= 14'h0949;
  filter_in_data[2578] <= 14'h3ecd;
  filter_in_data[2579] <= 14'h3920;
  filter_in_data[2580] <= 14'h0e6b;
  filter_in_data[2581] <= 14'h2b03;
  filter_in_data[2582] <= 14'h1a38;
  filter_in_data[2583] <= 14'h2226;
  filter_in_data[2584] <= 14'h1fbb;
  filter_in_data[2585] <= 14'h202e;
  filter_in_data[2586] <= 14'h1e2e;
  filter_in_data[2587] <= 14'h250a;
  filter_in_data[2588] <= 14'h1665;
  filter_in_data[2589] <= 14'h2f3e;
  filter_in_data[2590] <= 14'h0a62;
  filter_in_data[2591] <= 14'h3c68;
  filter_in_data[2592] <= 14'h3cbc;
  filter_in_data[2593] <= 14'h09e3;
  filter_in_data[2594] <= 14'h3005;
  filter_in_data[2595] <= 14'h154f;
  filter_in_data[2596] <= 14'h2652;
  filter_in_data[2597] <= 14'h1cf5;
  filter_in_data[2598] <= 14'h20f0;
  filter_in_data[2599] <= 14'h1ff6;
  filter_in_data[2600] <= 14'h2052;
  filter_in_data[2601] <= 14'h1e48;
  filter_in_data[2602] <= 14'h2423;
  filter_in_data[2603] <= 14'h1890;
  filter_in_data[2604] <= 14'h2b7a;
  filter_in_data[2605] <= 14'h0feb;
  filter_in_data[2606] <= 14'h3517;
  filter_in_data[2607] <= 14'h05ad;
  filter_in_data[2608] <= 14'h3fa1;
  filter_in_data[2609] <= 14'h3b28;
  filter_in_data[2610] <= 14'h09d8;
  filter_in_data[2611] <= 14'h3180;
  filter_in_data[2612] <= 14'h12b9;
  filter_in_data[2613] <= 14'h2993;
  filter_in_data[2614] <= 14'h198f;
  filter_in_data[2615] <= 14'h23eb;
  filter_in_data[2616] <= 14'h1dfa;
  filter_in_data[2617] <= 14'h20c2;
  filter_in_data[2618] <= 14'h1fe5;
  filter_in_data[2619] <= 14'h200b;
  filter_in_data[2620] <= 14'h1f78;
  filter_in_data[2621] <= 14'h2187;
  filter_in_data[2622] <= 14'h1d06;
  filter_in_data[2623] <= 14'h24d3;
  filter_in_data[2624] <= 14'h18fc;
  filter_in_data[2625] <= 14'h297c;
  filter_in_data[2626] <= 14'h13d2;
  filter_in_data[2627] <= 14'h2f0b;
  filter_in_data[2628] <= 14'h0dfa;
  filter_in_data[2629] <= 14'h3512;
  filter_in_data[2630] <= 14'h07dc;
  filter_in_data[2631] <= 14'h3b32;
  filter_in_data[2632] <= 14'h01cc;
  filter_in_data[2633] <= 14'h0120;
  filter_in_data[2634] <= 14'h3c0e;
  filter_in_data[2635] <= 14'h06a4;
  filter_in_data[2636] <= 14'h36ce;
  filter_in_data[2637] <= 14'h0b98;
  filter_in_data[2638] <= 14'h322a;
  filter_in_data[2639] <= 14'h0fea;
  filter_in_data[2640] <= 14'h2e2c;
  filter_in_data[2641] <= 14'h1393;
  filter_in_data[2642] <= 14'h2ad7;
  filter_in_data[2643] <= 14'h0000;
  filter_in_data[2644] <= 14'h0000;
  filter_in_data[2645] <= 14'h0000;
  filter_in_data[2646] <= 14'h0000;
  filter_in_data[2647] <= 14'h0000;
  filter_in_data[2648] <= 14'h0000;
  filter_in_data[2649] <= 14'h0000;
  filter_in_data[2650] <= 14'h0000;
  filter_in_data[2651] <= 14'h0000;
  filter_in_data[2652] <= 14'h0000;
  filter_in_data[2653] <= 14'h0000;
  filter_in_data[2654] <= 14'h0000;
  filter_in_data[2655] <= 14'h0000;
  filter_in_data[2656] <= 14'h0000;
  filter_in_data[2657] <= 14'h0000;
  filter_in_data[2658] <= 14'h0000;
  filter_in_data[2659] <= 14'h0000;
  filter_in_data[2660] <= 14'h0000;
  filter_in_data[2661] <= 14'h0000;
  filter_in_data[2662] <= 14'h0000;
  filter_in_data[2663] <= 14'h0000;
  filter_in_data[2664] <= 14'h0000;
  filter_in_data[2665] <= 14'h0000;
  filter_in_data[2666] <= 14'h0000;
  filter_in_data[2667] <= 14'h0000;
  filter_in_data[2668] <= 14'h0000;
  filter_in_data[2669] <= 14'h0000;
  filter_in_data[2670] <= 14'h0000;
  filter_in_data[2671] <= 14'h0000;
  filter_in_data[2672] <= 14'h0000;
  filter_in_data[2673] <= 14'h0000;
  filter_in_data[2674] <= 14'h0000;
  filter_in_data[2675] <= 14'h0000;
  filter_in_data[2676] <= 14'h0000;
  filter_in_data[2677] <= 14'h0000;
  filter_in_data[2678] <= 14'h0000;
  filter_in_data[2679] <= 14'h0000;
  filter_in_data[2680] <= 14'h0000;
  filter_in_data[2681] <= 14'h0000;
  filter_in_data[2682] <= 14'h0000;
  filter_in_data[2683] <= 14'h0000;
  filter_in_data[2684] <= 14'h0000;
  filter_in_data[2685] <= 14'h0000;
  filter_in_data[2686] <= 14'h0000;
  filter_in_data[2687] <= 14'h0000;
  filter_in_data[2688] <= 14'h0000;
  filter_in_data[2689] <= 14'h0000;
  filter_in_data[2690] <= 14'h0000;
  filter_in_data[2691] <= 14'h0000;
  filter_in_data[2692] <= 14'h0000;
  filter_in_data[2693] <= 14'h0000;
  filter_in_data[2694] <= 14'h0000;
  filter_in_data[2695] <= 14'h0000;
  filter_in_data[2696] <= 14'h0000;
  filter_in_data[2697] <= 14'h0000;
  filter_in_data[2698] <= 14'h0000;
  filter_in_data[2699] <= 14'h0000;
  filter_in_data[2700] <= 14'h0000;
  filter_in_data[2701] <= 14'h0000;
  filter_in_data[2702] <= 14'h0000;
  filter_in_data[2703] <= 14'h0000;
  filter_in_data[2704] <= 14'h0000;
  filter_in_data[2705] <= 14'h0000;
  filter_in_data[2706] <= 14'h0000;
  filter_in_data[2707] <= 14'h0000;
  filter_in_data[2708] <= 14'h0000;
  filter_in_data[2709] <= 14'h0000;
  filter_in_data[2710] <= 14'h0000;
  filter_in_data[2711] <= 14'h0000;
  filter_in_data[2712] <= 14'h0000;
  filter_in_data[2713] <= 14'h0000;
  filter_in_data[2714] <= 14'h0000;
  filter_in_data[2715] <= 14'h0000;
  filter_in_data[2716] <= 14'h0000;
  filter_in_data[2717] <= 14'h0000;
  filter_in_data[2718] <= 14'h0000;
  filter_in_data[2719] <= 14'h0000;
  filter_in_data[2720] <= 14'h0000;
  filter_in_data[2721] <= 14'h0000;
  filter_in_data[2722] <= 14'h0000;
  filter_in_data[2723] <= 14'h0000;
  filter_in_data[2724] <= 14'h0000;
  filter_in_data[2725] <= 14'h0000;
  filter_in_data[2726] <= 14'h0000;
  filter_in_data[2727] <= 14'h0000;
  filter_in_data[2728] <= 14'h0000;
  filter_in_data[2729] <= 14'h0000;
  filter_in_data[2730] <= 14'h0000;
  filter_in_data[2731] <= 14'h0000;
  filter_in_data[2732] <= 14'h0000;
  filter_in_data[2733] <= 14'h0000;
  filter_in_data[2734] <= 14'h0000;
  filter_in_data[2735] <= 14'h0000;
  filter_in_data[2736] <= 14'h0000;
  filter_in_data[2737] <= 14'h0000;
  filter_in_data[2738] <= 14'h0000;
  filter_in_data[2739] <= 14'h0000;
  filter_in_data[2740] <= 14'h0000;
  filter_in_data[2741] <= 14'h0000;
  filter_in_data[2742] <= 14'h0000;
  filter_in_data[2743] <= 14'h0000;
  filter_in_data[2744] <= 14'h0000;
  filter_in_data[2745] <= 14'h0000;
  filter_in_data[2746] <= 14'h0000;
  filter_in_data[2747] <= 14'h0000;
  filter_in_data[2748] <= 14'h0000;
  filter_in_data[2749] <= 14'h0000;
  filter_in_data[2750] <= 14'h0000;
  filter_in_data[2751] <= 14'h0000;
  filter_in_data[2752] <= 14'h0000;
  filter_in_data[2753] <= 14'h0000;
  filter_in_data[2754] <= 14'h0000;
  filter_in_data[2755] <= 14'h0000;
  filter_in_data[2756] <= 14'h0000;
  filter_in_data[2757] <= 14'h0000;
  filter_in_data[2758] <= 14'h0000;
  filter_in_data[2759] <= 14'h0000;
  filter_in_data[2760] <= 14'h0000;
  filter_in_data[2761] <= 14'h0000;
  filter_in_data[2762] <= 14'h2ba4;
  filter_in_data[2763] <= 14'h113d;
  filter_in_data[2764] <= 14'h2499;
  filter_in_data[2765] <= 14'h1bc7;
  filter_in_data[2766] <= 14'h241a;
  filter_in_data[2767] <= 14'h0a2c;
  filter_in_data[2768] <= 14'h268b;
  filter_in_data[2769] <= 14'h3b6f;
  filter_in_data[2770] <= 14'h3fcd;
  filter_in_data[2771] <= 14'h1733;
  filter_in_data[2772] <= 14'h3ff4;
  filter_in_data[2773] <= 14'h3d66;
  filter_in_data[2774] <= 14'h2630;
  filter_in_data[2775] <= 14'h34bb;
  filter_in_data[2776] <= 14'h07a2;
  filter_in_data[2777] <= 14'h2a2d;
  filter_in_data[2778] <= 14'h191e;
  filter_in_data[2779] <= 14'h2110;
  filter_in_data[2780] <= 14'h2708;
  filter_in_data[2781] <= 14'h2b72;
  filter_in_data[2782] <= 14'h32dd;
  filter_in_data[2783] <= 14'h3d77;
  filter_in_data[2784] <= 14'h36fc;
  filter_in_data[2785] <= 14'h2911;
  filter_in_data[2786] <= 14'h27d2;
  filter_in_data[2787] <= 14'h3dee;
  filter_in_data[2788] <= 14'h056d;
  filter_in_data[2789] <= 14'h155e;
  filter_in_data[2790] <= 14'h396b;
  filter_in_data[2791] <= 14'h02cb;
  filter_in_data[2792] <= 14'h2d19;
  filter_in_data[2793] <= 14'h2d0d;
  filter_in_data[2794] <= 14'h0c4b;
  filter_in_data[2795] <= 14'h2755;
  filter_in_data[2796] <= 14'h256f;
  filter_in_data[2797] <= 14'h1a83;
  filter_in_data[2798] <= 14'h0e20;
  filter_in_data[2799] <= 14'h11f5;
  filter_in_data[2800] <= 14'h1641;
  filter_in_data[2801] <= 14'h3660;
  filter_in_data[2802] <= 14'h2f8b;
  filter_in_data[2803] <= 14'h17bd;
  filter_in_data[2804] <= 14'h1171;
  filter_in_data[2805] <= 14'h03fc;
  filter_in_data[2806] <= 14'h0284;
  filter_in_data[2807] <= 14'h197e;
  filter_in_data[2808] <= 14'h1cf6;
  filter_in_data[2809] <= 14'h060f;
  filter_in_data[2810] <= 14'h0866;
  filter_in_data[2811] <= 14'h0799;
  filter_in_data[2812] <= 14'h2cf9;
  filter_in_data[2813] <= 14'h01de;
  filter_in_data[2814] <= 14'h32ec;
  filter_in_data[2815] <= 14'h1bb1;
  filter_in_data[2816] <= 14'h22d3;
  filter_in_data[2817] <= 14'h0c44;
  filter_in_data[2818] <= 14'h04a2;
  filter_in_data[2819] <= 14'h2dbf;
  filter_in_data[2820] <= 14'h1d0b;
  filter_in_data[2821] <= 14'h3b83;
  filter_in_data[2822] <= 14'h33b8;
  filter_in_data[2823] <= 14'h351e;
  filter_in_data[2824] <= 14'h0c44;
  filter_in_data[2825] <= 14'h16c4;
  filter_in_data[2826] <= 14'h018a;
  filter_in_data[2827] <= 14'h04fc;
  filter_in_data[2828] <= 14'h2809;
  filter_in_data[2829] <= 14'h2e55;
  filter_in_data[2830] <= 14'h0ea2;
  filter_in_data[2831] <= 14'h1fb2;
  filter_in_data[2832] <= 14'h3cfd;
  filter_in_data[2833] <= 14'h0e88;
  filter_in_data[2834] <= 14'h07af;
  filter_in_data[2835] <= 14'h0406;
  filter_in_data[2836] <= 14'h1d23;
  filter_in_data[2837] <= 14'h3c7a;
  filter_in_data[2838] <= 14'h0555;
  filter_in_data[2839] <= 14'h3c9d;
  filter_in_data[2840] <= 14'h37f0;
  filter_in_data[2841] <= 14'h1548;
  filter_in_data[2842] <= 14'h0f54;
  filter_in_data[2843] <= 14'h191b;
  filter_in_data[2844] <= 14'h3268;
  filter_in_data[2845] <= 14'h26eb;
  filter_in_data[2846] <= 14'h14ab;
  filter_in_data[2847] <= 14'h3c44;
  filter_in_data[2848] <= 14'h06af;
  filter_in_data[2849] <= 14'h130a;
  filter_in_data[2850] <= 14'h30c7;
  filter_in_data[2851] <= 14'h1346;
  filter_in_data[2852] <= 14'h1271;
  filter_in_data[2853] <= 14'h273d;
  filter_in_data[2854] <= 14'h004a;
  filter_in_data[2855] <= 14'h21aa;
  filter_in_data[2856] <= 14'h1ccb;
  filter_in_data[2857] <= 14'h1dba;
  filter_in_data[2858] <= 14'h07cf;
  filter_in_data[2859] <= 14'h040f;
  filter_in_data[2860] <= 14'h23d9;
  filter_in_data[2861] <= 14'h1917;
  filter_in_data[2862] <= 14'h37a1;
  filter_in_data[2863] <= 14'h08ef;
  filter_in_data[2864] <= 14'h1ad4;
  filter_in_data[2865] <= 14'h04af;
  filter_in_data[2866] <= 14'h2848;
  filter_in_data[2867] <= 14'h2c99;
  filter_in_data[2868] <= 14'h2607;
  filter_in_data[2869] <= 14'h2518;
  filter_in_data[2870] <= 14'h1054;
  filter_in_data[2871] <= 14'h288f;
  filter_in_data[2872] <= 14'h16dd;
  filter_in_data[2873] <= 14'h22de;
  filter_in_data[2874] <= 14'h355f;
  filter_in_data[2875] <= 14'h3e8a;
  filter_in_data[2876] <= 14'h15ef;
  filter_in_data[2877] <= 14'h0404;
  filter_in_data[2878] <= 14'h22cc;
  filter_in_data[2879] <= 14'h248f;
  filter_in_data[2880] <= 14'h19a9;
  filter_in_data[2881] <= 14'h2491;
  filter_in_data[2882] <= 14'h1ddd;
  filter_in_data[2883] <= 14'h02fd;
  filter_in_data[2884] <= 14'h3e70;
  filter_in_data[2885] <= 14'h32ec;
  filter_in_data[2886] <= 14'h1bee;
  filter_in_data[2887] <= 14'h20b1;
  filter_in_data[2888] <= 14'h3497;
  filter_in_data[2889] <= 14'h292e;
  filter_in_data[2890] <= 14'h31bc;
  filter_in_data[2891] <= 14'h135c;
  filter_in_data[2892] <= 14'h1c6c;
  filter_in_data[2893] <= 14'h0404;
  filter_in_data[2894] <= 14'h0630;
  filter_in_data[2895] <= 14'h0c85;
  filter_in_data[2896] <= 14'h2213;
  filter_in_data[2897] <= 14'h27ab;
  filter_in_data[2898] <= 14'h1e51;
  filter_in_data[2899] <= 14'h1d28;
  filter_in_data[2900] <= 14'h033c;
  filter_in_data[2901] <= 14'h2182;
  filter_in_data[2902] <= 14'h2658;
  filter_in_data[2903] <= 14'h13d9;
  filter_in_data[2904] <= 14'h2cb7;
  filter_in_data[2905] <= 14'h11ca;
  filter_in_data[2906] <= 14'h11f8;
  filter_in_data[2907] <= 14'h0f39;
  filter_in_data[2908] <= 14'h15db;
  filter_in_data[2909] <= 14'h2171;
  filter_in_data[2910] <= 14'h01ba;
  filter_in_data[2911] <= 14'h0c52;
  filter_in_data[2912] <= 14'h1dcd;
  filter_in_data[2913] <= 14'h0c9d;
  filter_in_data[2914] <= 14'h1689;
  filter_in_data[2915] <= 14'h383f;
  filter_in_data[2916] <= 14'h2ba0;
  filter_in_data[2917] <= 14'h16b3;
  filter_in_data[2918] <= 14'h2219;
  filter_in_data[2919] <= 14'h2d4e;
  filter_in_data[2920] <= 14'h087f;
  filter_in_data[2921] <= 14'h103e;
  filter_in_data[2922] <= 14'h0504;
  filter_in_data[2923] <= 14'h12d5;
  filter_in_data[2924] <= 14'h33aa;
  filter_in_data[2925] <= 14'h08eb;
  filter_in_data[2926] <= 14'h3fbb;
  filter_in_data[2927] <= 14'h151b;
  filter_in_data[2928] <= 14'h208a;
  filter_in_data[2929] <= 14'h31cf;
  filter_in_data[2930] <= 14'h2bb0;
  filter_in_data[2931] <= 14'h1eed;
  filter_in_data[2932] <= 14'h391b;
  filter_in_data[2933] <= 14'h213a;
  filter_in_data[2934] <= 14'h0b24;
  filter_in_data[2935] <= 14'h3ea4;
  filter_in_data[2936] <= 14'h1af7;
  filter_in_data[2937] <= 14'h3aae;
  filter_in_data[2938] <= 14'h2f5a;
  filter_in_data[2939] <= 14'h016c;
  filter_in_data[2940] <= 14'h26eb;
  filter_in_data[2941] <= 14'h1f10;
  filter_in_data[2942] <= 14'h2d88;
  filter_in_data[2943] <= 14'h1a51;
  filter_in_data[2944] <= 14'h2f62;
  filter_in_data[2945] <= 14'h0cb0;
  filter_in_data[2946] <= 14'h1f06;
  filter_in_data[2947] <= 14'h0565;
  filter_in_data[2948] <= 14'h0d2d;
  filter_in_data[2949] <= 14'h2b47;
  filter_in_data[2950] <= 14'h3859;
  filter_in_data[2951] <= 14'h004b;
  filter_in_data[2952] <= 14'h2b02;
  filter_in_data[2953] <= 14'h2d97;
  filter_in_data[2954] <= 14'h3fa7;
  filter_in_data[2955] <= 14'h042a;
  filter_in_data[2956] <= 14'h3402;
  filter_in_data[2957] <= 14'h18fd;
  filter_in_data[2958] <= 14'h26ad;
  filter_in_data[2959] <= 14'h0372;
  filter_in_data[2960] <= 14'h29c4;
  filter_in_data[2961] <= 14'h2207;
  filter_in_data[2962] <= 14'h0f1d;
  filter_in_data[2963] <= 14'h03a2;
  filter_in_data[2964] <= 14'h09df;
  filter_in_data[2965] <= 14'h1fd6;
  filter_in_data[2966] <= 14'h3c01;
  filter_in_data[2967] <= 14'h0632;
  filter_in_data[2968] <= 14'h30d0;
  filter_in_data[2969] <= 14'h208a;
  filter_in_data[2970] <= 14'h111f;
  filter_in_data[2971] <= 14'h11b3;
  filter_in_data[2972] <= 14'h1aa5;
  filter_in_data[2973] <= 14'h004a;
  filter_in_data[2974] <= 14'h03eb;
  filter_in_data[2975] <= 14'h28d9;
  filter_in_data[2976] <= 14'h26fd;
  filter_in_data[2977] <= 14'h310b;
  filter_in_data[2978] <= 14'h3636;
  filter_in_data[2979] <= 14'h101f;
  filter_in_data[2980] <= 14'h3205;
  filter_in_data[2981] <= 14'h2dda;
  filter_in_data[2982] <= 14'h061f;
  filter_in_data[2983] <= 14'h31e5;
  filter_in_data[2984] <= 14'h09d5;
  filter_in_data[2985] <= 14'h08ea;
  filter_in_data[2986] <= 14'h067f;
  filter_in_data[2987] <= 14'h06a1;
  filter_in_data[2988] <= 14'h3cb0;
  filter_in_data[2989] <= 14'h1656;
  filter_in_data[2990] <= 14'h3acb;
  filter_in_data[2991] <= 14'h14c0;
  filter_in_data[2992] <= 14'h28e6;
  filter_in_data[2993] <= 14'h3085;
  filter_in_data[2994] <= 14'h3eb7;
  filter_in_data[2995] <= 14'h315f;
  filter_in_data[2996] <= 14'h0409;
  filter_in_data[2997] <= 14'h204d;
  filter_in_data[2998] <= 14'h083b;
  filter_in_data[2999] <= 14'h3c35;
  filter_in_data[3000] <= 14'h1706;
  filter_in_data[3001] <= 14'h1708;
  filter_in_data[3002] <= 14'h03b8;
  filter_in_data[3003] <= 14'h118d;
  filter_in_data[3004] <= 14'h2716;
  filter_in_data[3005] <= 14'h07d4;
  filter_in_data[3006] <= 14'h37a1;
  filter_in_data[3007] <= 14'h23a0;
  filter_in_data[3008] <= 14'h2376;
  filter_in_data[3009] <= 14'h1f05;
  filter_in_data[3010] <= 14'h3994;
  filter_in_data[3011] <= 14'h080c;
  filter_in_data[3012] <= 14'h2caa;
  filter_in_data[3013] <= 14'h0f27;
  filter_in_data[3014] <= 14'h2881;
  filter_in_data[3015] <= 14'h3c50;
  filter_in_data[3016] <= 14'h1bf3;
  filter_in_data[3017] <= 14'h367f;
  filter_in_data[3018] <= 14'h150b;
  filter_in_data[3019] <= 14'h2290;
  filter_in_data[3020] <= 14'h2192;
  filter_in_data[3021] <= 14'h27ae;
  filter_in_data[3022] <= 14'h203c;
  filter_in_data[3023] <= 14'h288e;
  filter_in_data[3024] <= 14'h1e00;
  filter_in_data[3025] <= 14'h3e87;
  filter_in_data[3026] <= 14'h2ace;
  filter_in_data[3027] <= 14'h2f5a;
  filter_in_data[3028] <= 14'h2f3e;
  filter_in_data[3029] <= 14'h24e9;
  filter_in_data[3030] <= 14'h2d41;
  filter_in_data[3031] <= 14'h186d;
  filter_in_data[3032] <= 14'h3672;
  filter_in_data[3033] <= 14'h04e5;
  filter_in_data[3034] <= 14'h03f8;
  filter_in_data[3035] <= 14'h1b2b;
  filter_in_data[3036] <= 14'h0033;
  filter_in_data[3037] <= 14'h0373;
  filter_in_data[3038] <= 14'h196e;
  filter_in_data[3039] <= 14'h07b6;
  filter_in_data[3040] <= 14'h2f64;
  filter_in_data[3041] <= 14'h3ca5;
  filter_in_data[3042] <= 14'h327c;
  filter_in_data[3043] <= 14'h04f2;
  filter_in_data[3044] <= 14'h3462;
  filter_in_data[3045] <= 14'h1dee;
  filter_in_data[3046] <= 14'h22b4;
  filter_in_data[3047] <= 14'h3e8e;
  filter_in_data[3048] <= 14'h08f8;
  filter_in_data[3049] <= 14'h02e5;
  filter_in_data[3050] <= 14'h0637;
  filter_in_data[3051] <= 14'h27fd;
  filter_in_data[3052] <= 14'h0be3;
  filter_in_data[3053] <= 14'h387b;
  filter_in_data[3054] <= 14'h1897;
  filter_in_data[3055] <= 14'h372f;
  filter_in_data[3056] <= 14'h13ee;
  filter_in_data[3057] <= 14'h379d;
  filter_in_data[3058] <= 14'h1180;
  filter_in_data[3059] <= 14'h0203;
  filter_in_data[3060] <= 14'h10f7;
  filter_in_data[3061] <= 14'h245e;
  filter_in_data[3062] <= 14'h044a;
  filter_in_data[3063] <= 14'h2180;
  filter_in_data[3064] <= 14'h363e;
  filter_in_data[3065] <= 14'h0180;
  filter_in_data[3066] <= 14'h12a0;
  filter_in_data[3067] <= 14'h0e09;
  filter_in_data[3068] <= 14'h0fed;
  filter_in_data[3069] <= 14'h2e74;
  filter_in_data[3070] <= 14'h2a1b;
  filter_in_data[3071] <= 14'h2f4a;
  filter_in_data[3072] <= 14'h23ae;
  filter_in_data[3073] <= 14'h1198;
  filter_in_data[3074] <= 14'h25be;
  filter_in_data[3075] <= 14'h01f9;
  filter_in_data[3076] <= 14'h0b73;
  filter_in_data[3077] <= 14'h3d1c;
  filter_in_data[3078] <= 14'h0c7d;
  filter_in_data[3079] <= 14'h1ac6;
  filter_in_data[3080] <= 14'h3179;
  filter_in_data[3081] <= 14'h2104;
  filter_in_data[3082] <= 14'h1843;
  filter_in_data[3083] <= 14'h197f;
  filter_in_data[3084] <= 14'h1f09;
  filter_in_data[3085] <= 14'h1b2f;
  filter_in_data[3086] <= 14'h1ce7;
  filter_in_data[3087] <= 14'h2990;
  filter_in_data[3088] <= 14'h148a;
  filter_in_data[3089] <= 14'h297d;
  filter_in_data[3090] <= 14'h0142;
  filter_in_data[3091] <= 14'h0392;
  filter_in_data[3092] <= 14'h1ecd;
  filter_in_data[3093] <= 14'h2da4;
  filter_in_data[3094] <= 14'h2de9;
  filter_in_data[3095] <= 14'h07cc;
  filter_in_data[3096] <= 14'h0b20;
  filter_in_data[3097] <= 14'h09ba;
  filter_in_data[3098] <= 14'h3099;
  filter_in_data[3099] <= 14'h1997;
  filter_in_data[3100] <= 14'h044c;
  filter_in_data[3101] <= 14'h2e32;
  filter_in_data[3102] <= 14'h039c;
  filter_in_data[3103] <= 14'h1729;
  filter_in_data[3104] <= 14'h373e;
  filter_in_data[3105] <= 14'h2906;
  filter_in_data[3106] <= 14'h2fc8;
  filter_in_data[3107] <= 14'h0bec;
  filter_in_data[3108] <= 14'h2478;
  filter_in_data[3109] <= 14'h1319;
  filter_in_data[3110] <= 14'h38de;
  filter_in_data[3111] <= 14'h3e7f;
  filter_in_data[3112] <= 14'h16b5;
  filter_in_data[3113] <= 14'h26c5;
  filter_in_data[3114] <= 14'h3f46;
  filter_in_data[3115] <= 14'h11bc;
  filter_in_data[3116] <= 14'h2302;
  filter_in_data[3117] <= 14'h0d98;
  filter_in_data[3118] <= 14'h2d09;
  filter_in_data[3119] <= 14'h2741;
  filter_in_data[3120] <= 14'h1285;
  filter_in_data[3121] <= 14'h358b;
  filter_in_data[3122] <= 14'h125b;
  filter_in_data[3123] <= 14'h21b1;
  filter_in_data[3124] <= 14'h3890;
  filter_in_data[3125] <= 14'h19c7;
  filter_in_data[3126] <= 14'h036f;
  filter_in_data[3127] <= 14'h14f7;
  filter_in_data[3128] <= 14'h126a;
  filter_in_data[3129] <= 14'h1928;
  filter_in_data[3130] <= 14'h01fa;
  filter_in_data[3131] <= 14'h055f;
  filter_in_data[3132] <= 14'h0d9f;
  filter_in_data[3133] <= 14'h17d1;
  filter_in_data[3134] <= 14'h2453;
  filter_in_data[3135] <= 14'h1766;
  filter_in_data[3136] <= 14'h2784;
  filter_in_data[3137] <= 14'h1ef4;
  filter_in_data[3138] <= 14'h13fd;
  filter_in_data[3139] <= 14'h1686;
  filter_in_data[3140] <= 14'h194f;
  filter_in_data[3141] <= 14'h33f4;
  filter_in_data[3142] <= 14'h3619;
  filter_in_data[3143] <= 14'h2b3b;
  filter_in_data[3144] <= 14'h0f37;
  filter_in_data[3145] <= 14'h025c;
  filter_in_data[3146] <= 14'h0b0b;
  filter_in_data[3147] <= 14'h36c3;
  filter_in_data[3148] <= 14'h2073;
  filter_in_data[3149] <= 14'h0b4b;
  filter_in_data[3150] <= 14'h26c9;
  filter_in_data[3151] <= 14'h0af4;
  filter_in_data[3152] <= 14'h3dc6;
  filter_in_data[3153] <= 14'h0a13;
  filter_in_data[3154] <= 14'h0c3a;
  filter_in_data[3155] <= 14'h0288;
  filter_in_data[3156] <= 14'h3fe8;
  filter_in_data[3157] <= 14'h14e3;
  filter_in_data[3158] <= 14'h2114;
  filter_in_data[3159] <= 14'h1829;
  filter_in_data[3160] <= 14'h1dc7;
  filter_in_data[3161] <= 14'h05ce;
  filter_in_data[3162] <= 14'h3c90;
  filter_in_data[3163] <= 14'h1ad7;
  filter_in_data[3164] <= 14'h3b8b;
  filter_in_data[3165] <= 14'h119e;
  filter_in_data[3166] <= 14'h2491;
  filter_in_data[3167] <= 14'h22af;
  filter_in_data[3168] <= 14'h20ee;
  filter_in_data[3169] <= 14'h0b71;
  filter_in_data[3170] <= 14'h3f4b;
  filter_in_data[3171] <= 14'h0091;
  filter_in_data[3172] <= 14'h2fd1;
  filter_in_data[3173] <= 14'h0e3e;
  filter_in_data[3174] <= 14'h1af4;
  filter_in_data[3175] <= 14'h3f09;
  filter_in_data[3176] <= 14'h1546;
  filter_in_data[3177] <= 14'h16d1;
  filter_in_data[3178] <= 14'h3200;
  filter_in_data[3179] <= 14'h3b48;
  filter_in_data[3180] <= 14'h2183;
  filter_in_data[3181] <= 14'h2be3;
  filter_in_data[3182] <= 14'h0191;
  filter_in_data[3183] <= 14'h1302;
  filter_in_data[3184] <= 14'h2451;
  filter_in_data[3185] <= 14'h3ac6;
  filter_in_data[3186] <= 14'h0d9a;
  filter_in_data[3187] <= 14'h24ec;
  filter_in_data[3188] <= 14'h054b;
  filter_in_data[3189] <= 14'h1764;
  filter_in_data[3190] <= 14'h0b29;
  filter_in_data[3191] <= 14'h19de;
  filter_in_data[3192] <= 14'h08ac;
  filter_in_data[3193] <= 14'h30ef;
  filter_in_data[3194] <= 14'h2512;
  filter_in_data[3195] <= 14'h2ee6;
  filter_in_data[3196] <= 14'h0b20;
  filter_in_data[3197] <= 14'h0e1a;
  filter_in_data[3198] <= 14'h19ed;
  filter_in_data[3199] <= 14'h0afb;
  filter_in_data[3200] <= 14'h3f81;
  filter_in_data[3201] <= 14'h240f;
  filter_in_data[3202] <= 14'h0adc;
  filter_in_data[3203] <= 14'h315f;
  filter_in_data[3204] <= 14'h350d;
  filter_in_data[3205] <= 14'h2599;
  filter_in_data[3206] <= 14'h146a;
  filter_in_data[3207] <= 14'h3266;
  filter_in_data[3208] <= 14'h1852;
  filter_in_data[3209] <= 14'h29a8;
  filter_in_data[3210] <= 14'h2d48;
  filter_in_data[3211] <= 14'h1007;
  filter_in_data[3212] <= 14'h363c;
  filter_in_data[3213] <= 14'h261d;
  filter_in_data[3214] <= 14'h3ba9;
  filter_in_data[3215] <= 14'h0778;
  filter_in_data[3216] <= 14'h24e5;
  filter_in_data[3217] <= 14'h2b8a;
  filter_in_data[3218] <= 14'h175d;
  filter_in_data[3219] <= 14'h12db;
  filter_in_data[3220] <= 14'h0754;
  filter_in_data[3221] <= 14'h17e4;
  filter_in_data[3222] <= 14'h1e90;
  filter_in_data[3223] <= 14'h042b;
  filter_in_data[3224] <= 14'h3867;
  filter_in_data[3225] <= 14'h0899;
  filter_in_data[3226] <= 14'h134f;
  filter_in_data[3227] <= 14'h16b5;
  filter_in_data[3228] <= 14'h0ac0;
  filter_in_data[3229] <= 14'h1431;
  filter_in_data[3230] <= 14'h015d;
  filter_in_data[3231] <= 14'h1324;
  filter_in_data[3232] <= 14'h05da;
  filter_in_data[3233] <= 14'h0830;
  filter_in_data[3234] <= 14'h295a;
  filter_in_data[3235] <= 14'h3055;
  filter_in_data[3236] <= 14'h2a8b;
  filter_in_data[3237] <= 14'h34d0;
  filter_in_data[3238] <= 14'h3a79;
  filter_in_data[3239] <= 14'h31a0;
  filter_in_data[3240] <= 14'h26d8;
  filter_in_data[3241] <= 14'h2d65;
  filter_in_data[3242] <= 14'h2795;
  filter_in_data[3243] <= 14'h1e37;
  filter_in_data[3244] <= 14'h3e6a;
  filter_in_data[3245] <= 14'h3ea7;
  filter_in_data[3246] <= 14'h1be6;
  filter_in_data[3247] <= 14'h0886;
  filter_in_data[3248] <= 14'h1334;
  filter_in_data[3249] <= 14'h37c1;
  filter_in_data[3250] <= 14'h39a1;
  filter_in_data[3251] <= 14'h2c99;
  filter_in_data[3252] <= 14'h3dcd;
  filter_in_data[3253] <= 14'h11ca;
  filter_in_data[3254] <= 14'h0043;
  filter_in_data[3255] <= 14'h3f0b;
  filter_in_data[3256] <= 14'h129e;
  filter_in_data[3257] <= 14'h2de7;
  filter_in_data[3258] <= 14'h362f;
  filter_in_data[3259] <= 14'h02bd;
  filter_in_data[3260] <= 14'h1973;
  filter_in_data[3261] <= 14'h0f13;
  filter_in_data[3262] <= 14'h0a85;
  filter_in_data[3263] <= 14'h0525;
  filter_in_data[3264] <= 14'h36e8;
  filter_in_data[3265] <= 14'h0fbb;
  filter_in_data[3266] <= 14'h24ff;
  filter_in_data[3267] <= 14'h3449;
  filter_in_data[3268] <= 14'h2d7c;
  filter_in_data[3269] <= 14'h20ae;
  filter_in_data[3270] <= 14'h30e2;
  filter_in_data[3271] <= 14'h00ed;
  filter_in_data[3272] <= 14'h1c11;
  filter_in_data[3273] <= 14'h342e;
  filter_in_data[3274] <= 14'h2bb1;
  filter_in_data[3275] <= 14'h009a;
  filter_in_data[3276] <= 14'h170f;
  filter_in_data[3277] <= 14'h2422;
  filter_in_data[3278] <= 14'h2208;
  filter_in_data[3279] <= 14'h3a3a;
  filter_in_data[3280] <= 14'h2b7a;
  filter_in_data[3281] <= 14'h330b;
  filter_in_data[3282] <= 14'h2ed8;
  filter_in_data[3283] <= 14'h31e8;
  filter_in_data[3284] <= 14'h1b8e;
  filter_in_data[3285] <= 14'h2d6f;
  filter_in_data[3286] <= 14'h36a6;
  filter_in_data[3287] <= 14'h185d;
  filter_in_data[3288] <= 14'h2595;
  filter_in_data[3289] <= 14'h09c1;
  filter_in_data[3290] <= 14'h37d0;
  filter_in_data[3291] <= 14'h3bf1;
  filter_in_data[3292] <= 14'h16e3;
  filter_in_data[3293] <= 14'h3aac;
  filter_in_data[3294] <= 14'h20fc;
  filter_in_data[3295] <= 14'h3fbf;
  filter_in_data[3296] <= 14'h2c72;
  filter_in_data[3297] <= 14'h161c;
  filter_in_data[3298] <= 14'h28ca;
  filter_in_data[3299] <= 14'h2565;
  filter_in_data[3300] <= 14'h25f6;
  filter_in_data[3301] <= 14'h0035;
  filter_in_data[3302] <= 14'h1787;
  filter_in_data[3303] <= 14'h0b2f;
  filter_in_data[3304] <= 14'h1238;
  filter_in_data[3305] <= 14'h13af;
  filter_in_data[3306] <= 14'h2e54;
  filter_in_data[3307] <= 14'h34bb;
  filter_in_data[3308] <= 14'h1ccf;
  filter_in_data[3309] <= 14'h38eb;
  filter_in_data[3310] <= 14'h088b;
  filter_in_data[3311] <= 14'h2e9b;
  filter_in_data[3312] <= 14'h3083;
  filter_in_data[3313] <= 14'h0b1d;
  filter_in_data[3314] <= 14'h1af2;
  filter_in_data[3315] <= 14'h0506;
  filter_in_data[3316] <= 14'h1e34;
  filter_in_data[3317] <= 14'h3b32;
  filter_in_data[3318] <= 14'h2fbc;
  filter_in_data[3319] <= 14'h2987;
  filter_in_data[3320] <= 14'h280c;
  filter_in_data[3321] <= 14'h2abd;
  filter_in_data[3322] <= 14'h093b;
  filter_in_data[3323] <= 14'h165a;
  filter_in_data[3324] <= 14'h335f;
  filter_in_data[3325] <= 14'h3013;
  filter_in_data[3326] <= 14'h2983;
  filter_in_data[3327] <= 14'h101f;
  filter_in_data[3328] <= 14'h1670;
  filter_in_data[3329] <= 14'h231d;
  filter_in_data[3330] <= 14'h3515;
  filter_in_data[3331] <= 14'h01f5;
  filter_in_data[3332] <= 14'h12db;
  filter_in_data[3333] <= 14'h21c9;
  filter_in_data[3334] <= 14'h3d3d;
  filter_in_data[3335] <= 14'h1222;
  filter_in_data[3336] <= 14'h159e;
  filter_in_data[3337] <= 14'h2deb;
  filter_in_data[3338] <= 14'h0f69;
  filter_in_data[3339] <= 14'h3d83;
  filter_in_data[3340] <= 14'h22f9;
  filter_in_data[3341] <= 14'h35e0;
  filter_in_data[3342] <= 14'h24ad;
  filter_in_data[3343] <= 14'h11d9;
  filter_in_data[3344] <= 14'h31f2;
  filter_in_data[3345] <= 14'h10a3;
  filter_in_data[3346] <= 14'h20f0;
  filter_in_data[3347] <= 14'h2a16;
  filter_in_data[3348] <= 14'h299e;
  filter_in_data[3349] <= 14'h061e;
  filter_in_data[3350] <= 14'h1cac;
  filter_in_data[3351] <= 14'h0471;
  filter_in_data[3352] <= 14'h3f9f;
  filter_in_data[3353] <= 14'h1871;
  filter_in_data[3354] <= 14'h244d;
  filter_in_data[3355] <= 14'h144e;
  filter_in_data[3356] <= 14'h0f8f;
  filter_in_data[3357] <= 14'h1585;
  filter_in_data[3358] <= 14'h092a;
  filter_in_data[3359] <= 14'h3c12;
  filter_in_data[3360] <= 14'h12c9;
  filter_in_data[3361] <= 14'h08ea;
  filter_in_data[3362] <= 14'h00d5;
  filter_in_data[3363] <= 14'h24c9;
  filter_in_data[3364] <= 14'h2a4a;
  filter_in_data[3365] <= 14'h25f2;
  filter_in_data[3366] <= 14'h0c48;
  filter_in_data[3367] <= 14'h15a1;
  filter_in_data[3368] <= 14'h147e;
  filter_in_data[3369] <= 14'h27d6;
  filter_in_data[3370] <= 14'h1532;
  filter_in_data[3371] <= 14'h0a09;
  filter_in_data[3372] <= 14'h3101;
  filter_in_data[3373] <= 14'h209a;
  filter_in_data[3374] <= 14'h09f3;
  filter_in_data[3375] <= 14'h2234;
  filter_in_data[3376] <= 14'h05f7;
  filter_in_data[3377] <= 14'h1b25;
  filter_in_data[3378] <= 14'h350c;
  filter_in_data[3379] <= 14'h2693;
  filter_in_data[3380] <= 14'h1846;
  filter_in_data[3381] <= 14'h1bd7;
  filter_in_data[3382] <= 14'h1b08;
  filter_in_data[3383] <= 14'h219a;
  filter_in_data[3384] <= 14'h0f6e;
  filter_in_data[3385] <= 14'h1d4f;
  filter_in_data[3386] <= 14'h36d5;
  filter_in_data[3387] <= 14'h309f;
  filter_in_data[3388] <= 14'h0a46;
  filter_in_data[3389] <= 14'h3df4;
  filter_in_data[3390] <= 14'h381d;
  filter_in_data[3391] <= 14'h2ce4;
  filter_in_data[3392] <= 14'h36b6;
  filter_in_data[3393] <= 14'h34ee;
  filter_in_data[3394] <= 14'h1ca2;
  filter_in_data[3395] <= 14'h130d;
  filter_in_data[3396] <= 14'h2bf8;
  filter_in_data[3397] <= 14'h173c;
  filter_in_data[3398] <= 14'h3d5b;
  filter_in_data[3399] <= 14'h1bb9;
  filter_in_data[3400] <= 14'h3a31;
  filter_in_data[3401] <= 14'h35b6;
  filter_in_data[3402] <= 14'h2d68;
  filter_in_data[3403] <= 14'h04cd;
  filter_in_data[3404] <= 14'h2374;
  filter_in_data[3405] <= 14'h2dde;
  filter_in_data[3406] <= 14'h3a37;
  filter_in_data[3407] <= 14'h0a55;
  filter_in_data[3408] <= 14'h0b1f;
  filter_in_data[3409] <= 14'h0ec7;
  filter_in_data[3410] <= 14'h3a24;
  filter_in_data[3411] <= 14'h2637;
  filter_in_data[3412] <= 14'h1e3d;
  filter_in_data[3413] <= 14'h0a8b;
  filter_in_data[3414] <= 14'h0ed9;
  filter_in_data[3415] <= 14'h38b7;
  filter_in_data[3416] <= 14'h207c;
  filter_in_data[3417] <= 14'h3ebf;
  filter_in_data[3418] <= 14'h2fc1;
  filter_in_data[3419] <= 14'h198b;
  filter_in_data[3420] <= 14'h2509;
  filter_in_data[3421] <= 14'h0bc8;
  filter_in_data[3422] <= 14'h2809;
  filter_in_data[3423] <= 14'h2449;
  filter_in_data[3424] <= 14'h0586;
  filter_in_data[3425] <= 14'h1eff;
  filter_in_data[3426] <= 14'h2e33;
  filter_in_data[3427] <= 14'h3837;
  filter_in_data[3428] <= 14'h3e41;
  filter_in_data[3429] <= 14'h1990;
  filter_in_data[3430] <= 14'h208a;
  filter_in_data[3431] <= 14'h3340;
  filter_in_data[3432] <= 14'h0089;
  filter_in_data[3433] <= 14'h331a;
  filter_in_data[3434] <= 14'h08d1;
  filter_in_data[3435] <= 14'h043e;
  filter_in_data[3436] <= 14'h0f50;
  filter_in_data[3437] <= 14'h23f6;
  filter_in_data[3438] <= 14'h35f9;
  filter_in_data[3439] <= 14'h20ea;
  filter_in_data[3440] <= 14'h3127;
  filter_in_data[3441] <= 14'h10e5;
  filter_in_data[3442] <= 14'h050c;
  filter_in_data[3443] <= 14'h1b55;
  filter_in_data[3444] <= 14'h30b9;
  filter_in_data[3445] <= 14'h0b3f;
  filter_in_data[3446] <= 14'h0ff1;
  filter_in_data[3447] <= 14'h3054;
  filter_in_data[3448] <= 14'h3624;
  filter_in_data[3449] <= 14'h2a61;
  filter_in_data[3450] <= 14'h10eb;
  filter_in_data[3451] <= 14'h3f87;
  filter_in_data[3452] <= 14'h0985;
  filter_in_data[3453] <= 14'h0f19;
  filter_in_data[3454] <= 14'h0445;
  filter_in_data[3455] <= 14'h3106;
  filter_in_data[3456] <= 14'h05ef;
  filter_in_data[3457] <= 14'h0753;
  filter_in_data[3458] <= 14'h3db2;
  filter_in_data[3459] <= 14'h3ebb;
  filter_in_data[3460] <= 14'h0cc0;
  filter_in_data[3461] <= 14'h1368;
  filter_in_data[3462] <= 14'h3fb7;
  filter_in_data[3463] <= 14'h2b29;
  filter_in_data[3464] <= 14'h1801;
  filter_in_data[3465] <= 14'h2a4c;
  filter_in_data[3466] <= 14'h1758;
  filter_in_data[3467] <= 14'h2745;
  filter_in_data[3468] <= 14'h1186;
  filter_in_data[3469] <= 14'h2be0;
  filter_in_data[3470] <= 14'h28cd;
  filter_in_data[3471] <= 14'h3536;
  filter_in_data[3472] <= 14'h0a3c;
  filter_in_data[3473] <= 14'h315b;
  filter_in_data[3474] <= 14'h01dc;
  filter_in_data[3475] <= 14'h3463;
  filter_in_data[3476] <= 14'h2ec8;
  filter_in_data[3477] <= 14'h1adf;
  filter_in_data[3478] <= 14'h02e6;
  filter_in_data[3479] <= 14'h392a;
  filter_in_data[3480] <= 14'h12ab;
  filter_in_data[3481] <= 14'h02d7;
  filter_in_data[3482] <= 14'h1ffb;
  filter_in_data[3483] <= 14'h3270;
  filter_in_data[3484] <= 14'h181b;
  filter_in_data[3485] <= 14'h1bdc;
  filter_in_data[3486] <= 14'h16b2;
  filter_in_data[3487] <= 14'h3137;
  filter_in_data[3488] <= 14'h3aba;
  filter_in_data[3489] <= 14'h1a8b;
  filter_in_data[3490] <= 14'h26e5;
  filter_in_data[3491] <= 14'h162b;
  filter_in_data[3492] <= 14'h0ff2;
  filter_in_data[3493] <= 14'h063a;
  filter_in_data[3494] <= 14'h363c;
  filter_in_data[3495] <= 14'h04a3;
  filter_in_data[3496] <= 14'h389d;
  filter_in_data[3497] <= 14'h3859;
  filter_in_data[3498] <= 14'h3ce3;
  filter_in_data[3499] <= 14'h1605;
  filter_in_data[3500] <= 14'h04f7;
  filter_in_data[3501] <= 14'h327c;
  filter_in_data[3502] <= 14'h3c04;
  filter_in_data[3503] <= 14'h06fb;
  filter_in_data[3504] <= 14'h0e28;
  filter_in_data[3505] <= 14'h3b88;
  filter_in_data[3506] <= 14'h1994;
  filter_in_data[3507] <= 14'h1040;
  filter_in_data[3508] <= 14'h38b0;
  filter_in_data[3509] <= 14'h1c4d;
  filter_in_data[3510] <= 14'h2029;
  filter_in_data[3511] <= 14'h3626;
  filter_in_data[3512] <= 14'h0d0c;
  filter_in_data[3513] <= 14'h1a5c;
  filter_in_data[3514] <= 14'h1446;
  filter_in_data[3515] <= 14'h1944;
  filter_in_data[3516] <= 14'h2395;
  filter_in_data[3517] <= 14'h0f3f;
  filter_in_data[3518] <= 14'h3844;
  filter_in_data[3519] <= 14'h2269;
  filter_in_data[3520] <= 14'h2ed2;
  filter_in_data[3521] <= 14'h1b15;
  filter_in_data[3522] <= 14'h33eb;
  filter_in_data[3523] <= 14'h18cb;
  filter_in_data[3524] <= 14'h3261;
  filter_in_data[3525] <= 14'h30c4;
  filter_in_data[3526] <= 14'h0b89;
  filter_in_data[3527] <= 14'h123f;
  filter_in_data[3528] <= 14'h220c;
  filter_in_data[3529] <= 14'h2be4;
  filter_in_data[3530] <= 14'h3bcc;
  filter_in_data[3531] <= 14'h036a;
  filter_in_data[3532] <= 14'h2388;
  filter_in_data[3533] <= 14'h320f;
  filter_in_data[3534] <= 14'h0fc9;
  filter_in_data[3535] <= 14'h1f2f;
  filter_in_data[3536] <= 14'h2ea8;
  filter_in_data[3537] <= 14'h0f06;
  filter_in_data[3538] <= 14'h18e3;
  filter_in_data[3539] <= 14'h3ca0;
  filter_in_data[3540] <= 14'h2f7f;
  filter_in_data[3541] <= 14'h3b8a;
  filter_in_data[3542] <= 14'h3be7;
  filter_in_data[3543] <= 14'h3a3c;
  filter_in_data[3544] <= 14'h3954;
  filter_in_data[3545] <= 14'h3af3;
  filter_in_data[3546] <= 14'h0d7d;
  filter_in_data[3547] <= 14'h009b;
  filter_in_data[3548] <= 14'h0f3b;
  filter_in_data[3549] <= 14'h03d1;
  filter_in_data[3550] <= 14'h1916;
  filter_in_data[3551] <= 14'h019a;
  filter_in_data[3552] <= 14'h3431;
  filter_in_data[3553] <= 14'h104e;
  filter_in_data[3554] <= 14'h0e06;
  filter_in_data[3555] <= 14'h21b2;
  filter_in_data[3556] <= 14'h3f1d;
  filter_in_data[3557] <= 14'h2c62;
  filter_in_data[3558] <= 14'h0a8e;
  filter_in_data[3559] <= 14'h301b;
  filter_in_data[3560] <= 14'h023b;
  filter_in_data[3561] <= 14'h2266;
  filter_in_data[3562] <= 14'h0e52;
  filter_in_data[3563] <= 14'h164b;
  filter_in_data[3564] <= 14'h2e18;
  filter_in_data[3565] <= 14'h1829;
  filter_in_data[3566] <= 14'h1444;
  filter_in_data[3567] <= 14'h2c3c;
  filter_in_data[3568] <= 14'h1188;
  filter_in_data[3569] <= 14'h127f;
  filter_in_data[3570] <= 14'h0194;
  filter_in_data[3571] <= 14'h3ab4;
  filter_in_data[3572] <= 14'h1b0b;
  filter_in_data[3573] <= 14'h277e;
  filter_in_data[3574] <= 14'h1ab4;
  filter_in_data[3575] <= 14'h35bb;
  filter_in_data[3576] <= 14'h187e;
  filter_in_data[3577] <= 14'h1bba;
  filter_in_data[3578] <= 14'h2766;
  filter_in_data[3579] <= 14'h1385;
  filter_in_data[3580] <= 14'h25cc;
  filter_in_data[3581] <= 14'h1ee3;
  filter_in_data[3582] <= 14'h291d;
  filter_in_data[3583] <= 14'h2c50;
  filter_in_data[3584] <= 14'h0f14;
  filter_in_data[3585] <= 14'h06c9;
  filter_in_data[3586] <= 14'h10aa;
  filter_in_data[3587] <= 14'h397a;
  filter_in_data[3588] <= 14'h28de;
  filter_in_data[3589] <= 14'h06c6;
  filter_in_data[3590] <= 14'h3226;
  filter_in_data[3591] <= 14'h379c;
  filter_in_data[3592] <= 14'h1f14;
  filter_in_data[3593] <= 14'h2ad5;
  filter_in_data[3594] <= 14'h071f;
  filter_in_data[3595] <= 14'h1d41;
  filter_in_data[3596] <= 14'h15fa;
  filter_in_data[3597] <= 14'h30c3;
  filter_in_data[3598] <= 14'h22fd;
  filter_in_data[3599] <= 14'h06de;
  filter_in_data[3600] <= 14'h2aa0;
  filter_in_data[3601] <= 14'h23f8;
  filter_in_data[3602] <= 14'h132b;
  filter_in_data[3603] <= 14'h0475;
  filter_in_data[3604] <= 14'h3dd5;
  filter_in_data[3605] <= 14'h376d;
  filter_in_data[3606] <= 14'h310d;
  filter_in_data[3607] <= 14'h03a5;
  filter_in_data[3608] <= 14'h0a21;
  filter_in_data[3609] <= 14'h17c4;
  filter_in_data[3610] <= 14'h31ca;
  filter_in_data[3611] <= 14'h3a7b;
  filter_in_data[3612] <= 14'h3937;
  filter_in_data[3613] <= 14'h31a5;
  filter_in_data[3614] <= 14'h17a2;
  filter_in_data[3615] <= 14'h3c45;
  filter_in_data[3616] <= 14'h2f46;
  filter_in_data[3617] <= 14'h3881;
  filter_in_data[3618] <= 14'h0a91;
  filter_in_data[3619] <= 14'h208a;
  filter_in_data[3620] <= 14'h189d;
  filter_in_data[3621] <= 14'h04f4;
  filter_in_data[3622] <= 14'h0d77;
  filter_in_data[3623] <= 14'h35a2;
  filter_in_data[3624] <= 14'h1c5f;
  filter_in_data[3625] <= 14'h364e;
  filter_in_data[3626] <= 14'h0bda;
  filter_in_data[3627] <= 14'h3292;
  filter_in_data[3628] <= 14'h0a22;
  filter_in_data[3629] <= 14'h3a1a;
  filter_in_data[3630] <= 14'h129a;
  filter_in_data[3631] <= 14'h21d1;
  filter_in_data[3632] <= 14'h10c2;
  filter_in_data[3633] <= 14'h2b83;
  filter_in_data[3634] <= 14'h2383;
  filter_in_data[3635] <= 14'h0fb3;
  filter_in_data[3636] <= 14'h0e34;
  filter_in_data[3637] <= 14'h1590;
  filter_in_data[3638] <= 14'h3d3f;
  filter_in_data[3639] <= 14'h00b0;
  filter_in_data[3640] <= 14'h2c6c;
  filter_in_data[3641] <= 14'h115f;
  filter_in_data[3642] <= 14'h2085;
  filter_in_data[3643] <= 14'h13f8;
  filter_in_data[3644] <= 14'h0fb7;
  filter_in_data[3645] <= 14'h10b0;
  filter_in_data[3646] <= 14'h2f59;
  filter_in_data[3647] <= 14'h086e;
  filter_in_data[3648] <= 14'h0150;
  filter_in_data[3649] <= 14'h393c;
  filter_in_data[3650] <= 14'h1fc2;
  filter_in_data[3651] <= 14'h1c4c;
  filter_in_data[3652] <= 14'h0ca4;
  filter_in_data[3653] <= 14'h1e0e;
  filter_in_data[3654] <= 14'h1d50;
  filter_in_data[3655] <= 14'h2370;
  filter_in_data[3656] <= 14'h1aeb;
  filter_in_data[3657] <= 14'h20fb;
  filter_in_data[3658] <= 14'h0bbb;
  filter_in_data[3659] <= 14'h235d;
  filter_in_data[3660] <= 14'h1526;
  filter_in_data[3661] <= 14'h11ce;
  filter_in_data[3662] <= 14'h2aca;
  filter_in_data[3663] <= 14'h00b2;
  filter_in_data[3664] <= 14'h018d;
  filter_in_data[3665] <= 14'h0f37;
  filter_in_data[3666] <= 14'h2cc8;
  filter_in_data[3667] <= 14'h1894;
  filter_in_data[3668] <= 14'h229f;
  filter_in_data[3669] <= 14'h29fb;
  filter_in_data[3670] <= 14'h3117;
  filter_in_data[3671] <= 14'h13b2;
  filter_in_data[3672] <= 14'h234e;
  filter_in_data[3673] <= 14'h3738;
  filter_in_data[3674] <= 14'h3b9c;
  filter_in_data[3675] <= 14'h1589;
  filter_in_data[3676] <= 14'h2929;
  filter_in_data[3677] <= 14'h3c07;
  filter_in_data[3678] <= 14'h09ec;
  filter_in_data[3679] <= 14'h0927;
  filter_in_data[3680] <= 14'h0425;
  filter_in_data[3681] <= 14'h0213;
  filter_in_data[3682] <= 14'h3887;
  filter_in_data[3683] <= 14'h370b;
  filter_in_data[3684] <= 14'h3709;
  filter_in_data[3685] <= 14'h0356;
  filter_in_data[3686] <= 14'h0204;
  filter_in_data[3687] <= 14'h250e;
  filter_in_data[3688] <= 14'h06b4;
  filter_in_data[3689] <= 14'h39c3;
  filter_in_data[3690] <= 14'h0cd1;
  filter_in_data[3691] <= 14'h3b7b;
  filter_in_data[3692] <= 14'h1958;
  filter_in_data[3693] <= 14'h20bf;
  filter_in_data[3694] <= 14'h1d1f;
  filter_in_data[3695] <= 14'h052d;
  filter_in_data[3696] <= 14'h0b3f;
  filter_in_data[3697] <= 14'h142d;
  filter_in_data[3698] <= 14'h21e7;
  filter_in_data[3699] <= 14'h273a;
  filter_in_data[3700] <= 14'h2259;
  filter_in_data[3701] <= 14'h052c;
  filter_in_data[3702] <= 14'h3936;
  filter_in_data[3703] <= 14'h1b28;
  filter_in_data[3704] <= 14'h0de3;
  filter_in_data[3705] <= 14'h29f5;
  filter_in_data[3706] <= 14'h0744;
  filter_in_data[3707] <= 14'h0250;
  filter_in_data[3708] <= 14'h0369;
  filter_in_data[3709] <= 14'h1c03;
  filter_in_data[3710] <= 14'h20e8;
  filter_in_data[3711] <= 14'h22af;
  filter_in_data[3712] <= 14'h39cd;
  filter_in_data[3713] <= 14'h1e11;
  filter_in_data[3714] <= 14'h0774;
  filter_in_data[3715] <= 14'h0cd9;
  filter_in_data[3716] <= 14'h3c23;
  filter_in_data[3717] <= 14'h1ca8;
  filter_in_data[3718] <= 14'h11bd;
  filter_in_data[3719] <= 14'h371e;
  filter_in_data[3720] <= 14'h06fd;
  filter_in_data[3721] <= 14'h2a09;
  filter_in_data[3722] <= 14'h2998;
  filter_in_data[3723] <= 14'h06b2;
  filter_in_data[3724] <= 14'h3dfe;
  filter_in_data[3725] <= 14'h3080;
  filter_in_data[3726] <= 14'h2ef8;
  filter_in_data[3727] <= 14'h0321;
  filter_in_data[3728] <= 14'h0e6c;
  filter_in_data[3729] <= 14'h0219;
  filter_in_data[3730] <= 14'h375c;
  filter_in_data[3731] <= 14'h0756;
  filter_in_data[3732] <= 14'h06fe;
  filter_in_data[3733] <= 14'h25d1;
  filter_in_data[3734] <= 14'h323a;
  filter_in_data[3735] <= 14'h2edc;
  filter_in_data[3736] <= 14'h3a3a;
  filter_in_data[3737] <= 14'h19e8;
  filter_in_data[3738] <= 14'h3338;
  filter_in_data[3739] <= 14'h32ad;
  filter_in_data[3740] <= 14'h0550;
  filter_in_data[3741] <= 14'h2c94;
  filter_in_data[3742] <= 14'h2974;
  filter_in_data[3743] <= 14'h0d7b;
  filter_in_data[3744] <= 14'h3899;
  filter_in_data[3745] <= 14'h0822;
  filter_in_data[3746] <= 14'h38c6;
  filter_in_data[3747] <= 14'h010b;
  filter_in_data[3748] <= 14'h3743;
  filter_in_data[3749] <= 14'h22c9;
  filter_in_data[3750] <= 14'h3129;
  filter_in_data[3751] <= 14'h2b7a;
  filter_in_data[3752] <= 14'h023c;
  filter_in_data[3753] <= 14'h28cd;
  filter_in_data[3754] <= 14'h3432;
  filter_in_data[3755] <= 14'h30da;
  filter_in_data[3756] <= 14'h3ac7;
  filter_in_data[3757] <= 14'h04af;
  filter_in_data[3758] <= 14'h1f74;
  filter_in_data[3759] <= 14'h2540;
  filter_in_data[3760] <= 14'h2681;
  filter_in_data[3761] <= 14'h07a8;
  filter_in_data[3762] <= 14'h2687;
  filter_in_data[3763] <= 14'h389b;
  filter_in_data[3764] <= 14'h1c89;
  filter_in_data[3765] <= 14'h1f57;
  filter_in_data[3766] <= 14'h0ac7;
  filter_in_data[3767] <= 14'h35ff;
  filter_in_data[3768] <= 14'h0907;
  filter_in_data[3769] <= 14'h3187;
  filter_in_data[3770] <= 14'h196e;
  filter_in_data[3771] <= 14'h323b;
  filter_in_data[3772] <= 14'h3f6c;
  filter_in_data[3773] <= 14'h3e63;
  filter_in_data[3774] <= 14'h0ff0;
  filter_in_data[3775] <= 14'h3c0b;
  filter_in_data[3776] <= 14'h0e0f;
  filter_in_data[3777] <= 14'h07e7;
  filter_in_data[3778] <= 14'h08f9;
  filter_in_data[3779] <= 14'h2aa0;
  filter_in_data[3780] <= 14'h3168;
  filter_in_data[3781] <= 14'h1380;
  filter_in_data[3782] <= 14'h2b91;
  filter_in_data[3783] <= 14'h2b3b;
  filter_in_data[3784] <= 14'h1ab5;
  filter_in_data[3785] <= 14'h0035;
  filter_in_data[3786] <= 14'h0000;
  filter_in_data[3787] <= 14'h0000;
  filter_in_data[3788] <= 14'h0000;
  filter_in_data[3789] <= 14'h0000;
  filter_in_data[3790] <= 14'h0000;
  filter_in_data[3791] <= 14'h0000;
  filter_in_data[3792] <= 14'h0000;
  filter_in_data[3793] <= 14'h0000;
  filter_in_data[3794] <= 14'h0000;
  filter_in_data[3795] <= 14'h0000;
  filter_in_data[3796] <= 14'h0000;
  filter_in_data[3797] <= 14'h0000;
  filter_in_data[3798] <= 14'h0000;
  filter_in_data[3799] <= 14'h0000;
  filter_in_data[3800] <= 14'h0000;
  filter_in_data[3801] <= 14'h0000;
  filter_in_data[3802] <= 14'h0000;
  filter_in_data[3803] <= 14'h0000;
  filter_in_data[3804] <= 14'h0000;
  filter_in_data[3805] <= 14'h0000;
  filter_in_data[3806] <= 14'h0000;
  filter_in_data[3807] <= 14'h0000;
  filter_in_data[3808] <= 14'h0000;
  filter_in_data[3809] <= 14'h0000;
  filter_in_data[3810] <= 14'h0000;
  filter_in_data[3811] <= 14'h0000;
  filter_in_data[3812] <= 14'h0000;
  filter_in_data[3813] <= 14'h0000;
  filter_in_data[3814] <= 14'h0000;
  filter_in_data[3815] <= 14'h0000;
  filter_in_data[3816] <= 14'h0000;
  filter_in_data[3817] <= 14'h0000;
  filter_in_data[3818] <= 14'h0000;
  filter_in_data[3819] <= 14'h0000;
  filter_in_data[3820] <= 14'h0000;
  filter_in_data[3821] <= 14'h0000;
  filter_in_data[3822] <= 14'h0000;
  filter_in_data[3823] <= 14'h0000;
  filter_in_data[3824] <= 14'h0000;
  filter_in_data[3825] <= 14'h0000;
  filter_in_data[3826] <= 14'h0000;
  filter_in_data[3827] <= 14'h0000;
  filter_in_data[3828] <= 14'h0000;
  filter_in_data[3829] <= 14'h0000;
  filter_in_data[3830] <= 14'h0000;
  filter_in_data[3831] <= 14'h0000;
  filter_in_data[3832] <= 14'h0000;
  filter_in_data[3833] <= 14'h0000;
  filter_in_data[3834] <= 14'h0000;
  filter_in_data[3835] <= 14'h0000;
  filter_in_data[3836] <= 14'h0000;
  filter_in_data[3837] <= 14'h0000;
  filter_in_data[3838] <= 14'h0000;
  filter_in_data[3839] <= 14'h0000;
  filter_in_data[3840] <= 14'h0000;
  filter_in_data[3841] <= 14'h0000;
  filter_in_data[3842] <= 14'h0000;
  filter_in_data[3843] <= 14'h0000;
  filter_in_data[3844] <= 14'h0000;
  filter_in_data[3845] <= 14'h0000;
  filter_in_data[3846] <= 14'h0000;
  filter_in_data[3847] <= 14'h0000;
  filter_in_data[3848] <= 14'h0000;
  filter_in_data[3849] <= 14'h0000;
  filter_in_data[3850] <= 14'h0000;
  filter_in_data[3851] <= 14'h0000;
  filter_in_data[3852] <= 14'h0000;
  filter_in_data[3853] <= 14'h0000;
  filter_in_data[3854] <= 14'h0000;
  filter_in_data[3855] <= 14'h0000;
  filter_in_data[3856] <= 14'h0000;
  filter_in_data[3857] <= 14'h0000;
  filter_in_data[3858] <= 14'h0000;
  filter_in_data[3859] <= 14'h0000;
  filter_in_data[3860] <= 14'h0000;
  filter_in_data[3861] <= 14'h0000;
  filter_in_data[3862] <= 14'h0000;
  filter_in_data[3863] <= 14'h0000;
  filter_in_data[3864] <= 14'h0000;
  filter_in_data[3865] <= 14'h0000;
  filter_in_data[3866] <= 14'h0000;
  filter_in_data[3867] <= 14'h0000;
  filter_in_data[3868] <= 14'h0000;
  filter_in_data[3869] <= 14'h0000;
  filter_in_data[3870] <= 14'h0000;
  filter_in_data[3871] <= 14'h0000;
  filter_in_data[3872] <= 14'h0000;
  filter_in_data[3873] <= 14'h0000;
  filter_in_data[3874] <= 14'h0000;
  filter_in_data[3875] <= 14'h0000;
  filter_in_data[3876] <= 14'h0000;
  filter_in_data[3877] <= 14'h0000;
  filter_in_data[3878] <= 14'h0000;
  filter_in_data[3879] <= 14'h0000;
  filter_in_data[3880] <= 14'h0000;
  filter_in_data[3881] <= 14'h0000;
  filter_in_data[3882] <= 14'h0000;
  filter_in_data[3883] <= 14'h0000;
  filter_in_data[3884] <= 14'h0000;
  filter_in_data[3885] <= 14'h0000;
  filter_in_data[3886] <= 14'h0000;
  filter_in_data[3887] <= 14'h0000;
  filter_in_data[3888] <= 14'h0000;
  filter_in_data[3889] <= 14'h0000;
  filter_in_data[3890] <= 14'h0000;
  filter_in_data[3891] <= 14'h0000;
  filter_in_data[3892] <= 14'h0000;
  filter_in_data[3893] <= 14'h0000;
  filter_in_data[3894] <= 14'h0000;
  filter_in_data[3895] <= 14'h0000;
  filter_in_data[3896] <= 14'h0000;
  filter_in_data[3897] <= 14'h0000;
  filter_in_data[3898] <= 14'h0000;
  filter_in_data[3899] <= 14'h0000;
  filter_in_data[3900] <= 14'h0000;
  filter_in_data[3901] <= 14'h0000;
  filter_in_data[3902] <= 14'h0000;
  filter_in_data[3903] <= 14'h0000;
  filter_in_data[3904] <= 14'h0000;


  @(negedge clock);
    reset = 0;
  @(negedge clock);
    reset = 1;
    clk_enable = 1;
  @(negedge clock);
    reset = 0;
    // next two lines below should be added    
    $set_toggle_region(filt);
    $toggle_start();
    for (int i = 0; i < 3905; i += 1) begin
      filt_in = filter_in_data[i];
      for (int j = 0; j < 60; j+=1) begin
          @(negedge clock);
      end
      $display("Loop: %d filt_in: %d filt_out[0]: %d ", i, filt_in, filt_out[0]);
    end
    
    // next two lines should be added
    $toggle_stop();
    $toggle_report("rand.saif", 1e-9, filt);
    $finish;
	end
endmodule
